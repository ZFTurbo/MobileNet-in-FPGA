module border(
    input clk, go,
    input [14:0] i,
    input [7:0] matrix,
    output reg [1:0] prov
);
	always @(posedge clk)
	begin	
		if (go == 1)
		begin
			prov = 0;
				if ((i == 1*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 2*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 3*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 4*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 5*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 6*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 7*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 8*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 9*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 10*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 11*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 12*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 13*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 14*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 15*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 16*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 17*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 18*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 19*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 20*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 21*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 22*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 23*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 24*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 25*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 26*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 27*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 28*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 29*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 30*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 31*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 32*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 33*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 34*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 35*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 36*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 37*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 38*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 39*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 40*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 41*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 42*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 43*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 44*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 45*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 46*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 47*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 48*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 49*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 50*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 51*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 52*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 53*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 54*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 55*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 56*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 57*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 58*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 59*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 60*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 61*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 62*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 63*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 64*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 65*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 66*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 67*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 68*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 69*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 70*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 71*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 72*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 73*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 74*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 75*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 76*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 77*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 78*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 79*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 80*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 81*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 82*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 83*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 84*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 85*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 86*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 87*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 88*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 89*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 90*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 91*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 92*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 93*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 94*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 95*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 96*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 97*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 98*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 99*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 100*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 101*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 102*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 103*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 104*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 105*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 106*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 107*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 108*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 109*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 110*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 111*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 112*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 113*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 114*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 115*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 116*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 117*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 118*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 119*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 120*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 121*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 122*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 123*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 124*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 125*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 126*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 127*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;
				if ((i == 128*matrix-1'b1) && (prov != 2'b10))	prov = 2'b10;

               if ((i == 0*matrix) && (prov != 2'b11))		    prov = 2'b11;
               if ((i == 1*matrix) && (prov != 2'b11))		    prov = 2'b11;
               if ((i == 2*matrix) && (prov != 2'b11))		    prov = 2'b11;
               if ((i == 3*matrix) && (prov != 2'b11))		    prov = 2'b11;
               if ((i == 4*matrix) && (prov != 2'b11))		    prov = 2'b11;
               if ((i == 5*matrix) && (prov != 2'b11))		    prov = 2'b11;
               if ((i == 6*matrix) && (prov != 2'b11))		    prov = 2'b11;
               if ((i == 7*matrix) && (prov != 2'b11))		    prov = 2'b11;
               if ((i == 8*matrix) && (prov != 2'b11))		    prov = 2'b11;
               if ((i == 9*matrix) && (prov != 2'b11))		    prov = 2'b11;
               if ((i == 10*matrix) && (prov != 2'b11))		    prov = 2'b11;
               if ((i == 11*matrix) && (prov != 2'b11))		    prov = 2'b11;
               if ((i == 12*matrix) && (prov != 2'b11))		    prov = 2'b11;
               if ((i == 13*matrix) && (prov != 2'b11))		    prov = 2'b11;
               if ((i == 14*matrix) && (prov != 2'b11))		    prov = 2'b11;
               if ((i == 15*matrix) && (prov != 2'b11))		    prov = 2'b11;
               if ((i == 16*matrix) && (prov != 2'b11))		    prov = 2'b11;
               if ((i == 17*matrix) && (prov != 2'b11))		    prov = 2'b11;
               if ((i == 18*matrix) && (prov != 2'b11))		    prov = 2'b11;
               if ((i == 19*matrix) && (prov != 2'b11))		    prov = 2'b11;
               if ((i == 20*matrix) && (prov != 2'b11))		    prov = 2'b11;
               if ((i == 21*matrix) && (prov != 2'b11))		    prov = 2'b11;
               if ((i == 22*matrix) && (prov != 2'b11))		    prov = 2'b11;
               if ((i == 23*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 24*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 25*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 26*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 27*matrix) && (prov != 2'b11))		    prov = 2'b11;
               if ((i == 28*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 29*matrix) && (prov != 2'b11))		    prov = 2'b11;
               if ((i == 30*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 31*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 32*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 33*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 34*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 35*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 36*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 37*matrix) && (prov != 2'b11))	        prov = 2'b11;
               if ((i == 38*matrix) && (prov != 2'b11))		    prov = 2'b11;
               if ((i == 39*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 40*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 41*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 42*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 43*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 44*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 45*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 46*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 47*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 48*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 49*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 50*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 51*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 52*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 53*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 54*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 55*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 56*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 57*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 58*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 59*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 60*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 61*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 62*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 63*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 64*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 65*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 66*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 67*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 68*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 69*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 70*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 71*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 72*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 73*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 74*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 75*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 76*matrix) && (prov != 2'b11))		    prov = 2'b11;
               if ((i == 77*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 78*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 79*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 80*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 81*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 82*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 83*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 84*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 85*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 86*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 87*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 88*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 89*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 90*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 91*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 92*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 93*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 94*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 95*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 96*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 97*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 98*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 99*matrix) && (prov != 2'b11))	    	prov = 2'b11;
               if ((i == 100*matrix) && (prov != 2'b11))	    prov = 2'b11;
               if ((i == 101*matrix) && (prov != 2'b11))		prov = 2'b11;
               if ((i == 102*matrix) && (prov != 2'b11))		prov = 2'b11;
               if ((i == 103*matrix) && (prov != 2'b11))		prov = 2'b11;
               if ((i == 104*matrix) && (prov != 2'b11))		prov = 2'b11;
               if ((i == 105*matrix) && (prov != 2'b11))		prov = 2'b11;
               if ((i == 106*matrix) && (prov != 2'b11))		prov = 2'b11;
               if ((i == 107*matrix) && (prov != 2'b11))		prov = 2'b11;
               if ((i == 108*matrix) && (prov != 2'b11))		prov = 2'b11;
               if ((i == 109*matrix) && (prov != 2'b11))		prov = 2'b11;
               if ((i == 110*matrix) && (prov != 2'b11))		prov = 2'b11;
               if ((i == 111*matrix) && (prov != 2'b11))		prov = 2'b11;
               if ((i == 112*matrix) && (prov != 2'b11))		prov = 2'b11;
               if ((i == 113*matrix) && (prov != 2'b11))		prov = 2'b11;
               if ((i == 114*matrix) && (prov != 2'b11))		prov = 2'b11;
               if ((i == 115*matrix) && (prov != 2'b11))		prov = 2'b11;
               if ((i == 116*matrix) && (prov != 2'b11))		prov = 2'b11;
               if ((i == 117*matrix) && (prov != 2'b11))		prov = 2'b11;
               if ((i == 118*matrix) && (prov != 2'b11))		prov = 2'b11;
               if ((i == 119*matrix) && (prov != 2'b11))		prov = 2'b11;
               if ((i == 120*matrix) && (prov != 2'b11))		prov = 2'b11;
               if ((i == 121*matrix) && (prov != 2'b11))		prov = 2'b11;
               if ((i == 122*matrix) && (prov != 2'b11))		prov = 2'b11;
               if ((i == 123*matrix) && (prov != 2'b11))		prov = 2'b11;
               if ((i == 124*matrix) && (prov != 2'b11))		prov = 2'b11;
               if ((i == 125*matrix) && (prov != 2'b11))		prov = 2'b11;
               if ((i == 126*matrix) && (prov != 2'b11))		prov = 2'b11;
               if ((i == 127*matrix) && (prov != 2'b11))		prov = 2'b11;
               if ((i == 128*matrix) && (prov != 2'b11))		prov = 2'b11;
		end
		else
			prov = 0;
	end
endmodule
