module scale_picture(
clk,
rst,
valid_data,
r,
g,
b,
x,
y,
r_out,
g_out,
b_out,
addr_out,
valid_data_out,
test
);
input clk,rst;
input valid_data;
input [7:0] r;
input [7:0] g;
input [7:0] b;
input [8:0] x,y;
output reg [7:0] r_out;
output reg [7:0] g_out;
output reg [7:0] b_out;
output [16:0] addr_out;
output reg valid_data_out;
output wire [15:0] test;

wire [16:0] addr_data;
reg [16:0] addr_k;
reg [16:0] i;

reg [7:0] data_mem_red [0:321];
reg [7:0] data_mem_green [0:321];
reg [7:0] data_mem_blue [0:321];

reg [7:0] p1_red,p2_red,p3_red,p4_red;
reg [7:0] p1_green,p2_green,p3_green,p4_green;
reg [7:0] p1_blue,p2_blue,p3_blue,p4_blue;

reg [23:0] r_res,g_res,b_res;

reg [7:0] razn_h_mem [0:128*128-1];
reg [7:0] razn_w_mem [0:128*128-1];
reg [15:0] k1,k2,k3,k4;

reg [16:0] mem_k_index [0:128*128-1];

always @(posedge clk or negedge rst)
	if (!rst) 
		begin
			addr_k = 0;
			k1 = 0;
			k2 = 0;
			k3 = 0;
			k4 = 0;
			r_out = 0;
			g_out = 0;
			b_out = 0;
			valid_data_out = 0;
		end
	else
		begin
		if (valid_data)
			begin
				data_mem_red[320+1] = r;
				data_mem_green[320+1] = g;
				data_mem_blue[320+1] = b;
				if ((addr_data+(320+1)) == ((y*320 + x)))
					begin
						valid_data_out = 1;

						k1 = (255 - razn_h_mem[addr_k]) * (255 - razn_w_mem[addr_k]);
						k2 = (255 - razn_h_mem[addr_k]) * razn_w_mem[addr_k];
						k3 = razn_h_mem[addr_k] * razn_w_mem[addr_k];
						k4 = razn_h_mem[addr_k] * (255 - razn_w_mem[addr_k]);
						
						p1_red = data_mem_red[0];
						p1_green = data_mem_green[0];
						p1_blue = data_mem_blue[0];
						
						p2_red = data_mem_red[320];
						p2_green = data_mem_green[320];
						p2_blue = data_mem_blue[320];
						
						p3_red = data_mem_red[321];
						p3_green = data_mem_green[321];
						p3_blue = data_mem_blue[321];
						
						p4_red = data_mem_red[1];
						p4_green = data_mem_green[1];
						p4_blue = data_mem_blue[1];
						
						r_res = p1_red * k1 + p2_red * k2 + p3_red * k3 + p4_red * k4;
						r_out = r_res[23:16];
						
						g_res = p1_green * k1 + p2_green * k2 + p3_green * k3 + p4_green * k4;
						g_out = g_res[23:16];
						
						b_res = p1_blue * k1 + p2_blue * k2 + p3_blue * k3 + p4_blue * k4;
						b_out = b_res[23:16];
						
						if (addr_k<128*128-1) addr_k = addr_k + 1;
						else addr_k = 0;
					end
				else valid_data_out = 0;
				for (i = 1; i <=321; i = i + 1)
					begin
						data_mem_red[i-1] = data_mem_red[i];
						data_mem_green[i-1] = data_mem_green[i];
						data_mem_blue[i-1] = data_mem_blue[i];
					end
			end
		else
			begin
				valid_data_out = 0;
			end
		end

assign test = addr_data[15:0];
assign addr_data = mem_k_index[addr_k];
assign addr_out = addr_k;
	
initial //mem_k_index
begin
mem_k_index[0] = 0;
mem_k_index[1] = 2;
mem_k_index[2] = 5;
mem_k_index[3] = 7;
mem_k_index[4] = 10;
mem_k_index[5] = 12;
mem_k_index[6] = 15;
mem_k_index[7] = 17;
mem_k_index[8] = 20;
mem_k_index[9] = 22;
mem_k_index[10] = 25;
mem_k_index[11] = 27;
mem_k_index[12] = 30;
mem_k_index[13] = 32;
mem_k_index[14] = 35;
mem_k_index[15] = 37;
mem_k_index[16] = 40;
mem_k_index[17] = 42;
mem_k_index[18] = 45;
mem_k_index[19] = 47;
mem_k_index[20] = 50;
mem_k_index[21] = 52;
mem_k_index[22] = 55;
mem_k_index[23] = 57;
mem_k_index[24] = 60;
mem_k_index[25] = 62;
mem_k_index[26] = 65;
mem_k_index[27] = 67;
mem_k_index[28] = 70;
mem_k_index[29] = 72;
mem_k_index[30] = 75;
mem_k_index[31] = 77;
mem_k_index[32] = 80;
mem_k_index[33] = 82;
mem_k_index[34] = 85;
mem_k_index[35] = 87;
mem_k_index[36] = 90;
mem_k_index[37] = 92;
mem_k_index[38] = 95;
mem_k_index[39] = 97;
mem_k_index[40] = 100;
mem_k_index[41] = 102;
mem_k_index[42] = 105;
mem_k_index[43] = 108;
mem_k_index[44] = 110;
mem_k_index[45] = 113;
mem_k_index[46] = 115;
mem_k_index[47] = 118;
mem_k_index[48] = 120;
mem_k_index[49] = 123;
mem_k_index[50] = 125;
mem_k_index[51] = 128;
mem_k_index[52] = 130;
mem_k_index[53] = 133;
mem_k_index[54] = 135;
mem_k_index[55] = 138;
mem_k_index[56] = 140;
mem_k_index[57] = 143;
mem_k_index[58] = 145;
mem_k_index[59] = 148;
mem_k_index[60] = 150;
mem_k_index[61] = 153;
mem_k_index[62] = 155;
mem_k_index[63] = 158;
mem_k_index[64] = 160;
mem_k_index[65] = 163;
mem_k_index[66] = 165;
mem_k_index[67] = 168;
mem_k_index[68] = 170;
mem_k_index[69] = 173;
mem_k_index[70] = 175;
mem_k_index[71] = 178;
mem_k_index[72] = 180;
mem_k_index[73] = 183;
mem_k_index[74] = 185;
mem_k_index[75] = 188;
mem_k_index[76] = 190;
mem_k_index[77] = 193;
mem_k_index[78] = 195;
mem_k_index[79] = 198;
mem_k_index[80] = 200;
mem_k_index[81] = 203;
mem_k_index[82] = 205;
mem_k_index[83] = 208;
mem_k_index[84] = 210;
mem_k_index[85] = 213;
mem_k_index[86] = 216;
mem_k_index[87] = 218;
mem_k_index[88] = 221;
mem_k_index[89] = 223;
mem_k_index[90] = 226;
mem_k_index[91] = 228;
mem_k_index[92] = 231;
mem_k_index[93] = 233;
mem_k_index[94] = 236;
mem_k_index[95] = 238;
mem_k_index[96] = 241;
mem_k_index[97] = 243;
mem_k_index[98] = 246;
mem_k_index[99] = 248;
mem_k_index[100] = 251;
mem_k_index[101] = 253;
mem_k_index[102] = 256;
mem_k_index[103] = 258;
mem_k_index[104] = 261;
mem_k_index[105] = 263;
mem_k_index[106] = 266;
mem_k_index[107] = 268;
mem_k_index[108] = 271;
mem_k_index[109] = 273;
mem_k_index[110] = 276;
mem_k_index[111] = 278;
mem_k_index[112] = 281;
mem_k_index[113] = 283;
mem_k_index[114] = 286;
mem_k_index[115] = 288;
mem_k_index[116] = 291;
mem_k_index[117] = 293;
mem_k_index[118] = 296;
mem_k_index[119] = 298;
mem_k_index[120] = 301;
mem_k_index[121] = 303;
mem_k_index[122] = 306;
mem_k_index[123] = 308;
mem_k_index[124] = 311;
mem_k_index[125] = 313;
mem_k_index[126] = 316;
mem_k_index[127] = 318;
mem_k_index[128] = 320;
mem_k_index[129] = 322;
mem_k_index[130] = 325;
mem_k_index[131] = 327;
mem_k_index[132] = 330;
mem_k_index[133] = 332;
mem_k_index[134] = 335;
mem_k_index[135] = 337;
mem_k_index[136] = 340;
mem_k_index[137] = 342;
mem_k_index[138] = 345;
mem_k_index[139] = 347;
mem_k_index[140] = 350;
mem_k_index[141] = 352;
mem_k_index[142] = 355;
mem_k_index[143] = 357;
mem_k_index[144] = 360;
mem_k_index[145] = 362;
mem_k_index[146] = 365;
mem_k_index[147] = 367;
mem_k_index[148] = 370;
mem_k_index[149] = 372;
mem_k_index[150] = 375;
mem_k_index[151] = 377;
mem_k_index[152] = 380;
mem_k_index[153] = 382;
mem_k_index[154] = 385;
mem_k_index[155] = 387;
mem_k_index[156] = 390;
mem_k_index[157] = 392;
mem_k_index[158] = 395;
mem_k_index[159] = 397;
mem_k_index[160] = 400;
mem_k_index[161] = 402;
mem_k_index[162] = 405;
mem_k_index[163] = 407;
mem_k_index[164] = 410;
mem_k_index[165] = 412;
mem_k_index[166] = 415;
mem_k_index[167] = 417;
mem_k_index[168] = 420;
mem_k_index[169] = 422;
mem_k_index[170] = 425;
mem_k_index[171] = 428;
mem_k_index[172] = 430;
mem_k_index[173] = 433;
mem_k_index[174] = 435;
mem_k_index[175] = 438;
mem_k_index[176] = 440;
mem_k_index[177] = 443;
mem_k_index[178] = 445;
mem_k_index[179] = 448;
mem_k_index[180] = 450;
mem_k_index[181] = 453;
mem_k_index[182] = 455;
mem_k_index[183] = 458;
mem_k_index[184] = 460;
mem_k_index[185] = 463;
mem_k_index[186] = 465;
mem_k_index[187] = 468;
mem_k_index[188] = 470;
mem_k_index[189] = 473;
mem_k_index[190] = 475;
mem_k_index[191] = 478;
mem_k_index[192] = 480;
mem_k_index[193] = 483;
mem_k_index[194] = 485;
mem_k_index[195] = 488;
mem_k_index[196] = 490;
mem_k_index[197] = 493;
mem_k_index[198] = 495;
mem_k_index[199] = 498;
mem_k_index[200] = 500;
mem_k_index[201] = 503;
mem_k_index[202] = 505;
mem_k_index[203] = 508;
mem_k_index[204] = 510;
mem_k_index[205] = 513;
mem_k_index[206] = 515;
mem_k_index[207] = 518;
mem_k_index[208] = 520;
mem_k_index[209] = 523;
mem_k_index[210] = 525;
mem_k_index[211] = 528;
mem_k_index[212] = 530;
mem_k_index[213] = 533;
mem_k_index[214] = 536;
mem_k_index[215] = 538;
mem_k_index[216] = 541;
mem_k_index[217] = 543;
mem_k_index[218] = 546;
mem_k_index[219] = 548;
mem_k_index[220] = 551;
mem_k_index[221] = 553;
mem_k_index[222] = 556;
mem_k_index[223] = 558;
mem_k_index[224] = 561;
mem_k_index[225] = 563;
mem_k_index[226] = 566;
mem_k_index[227] = 568;
mem_k_index[228] = 571;
mem_k_index[229] = 573;
mem_k_index[230] = 576;
mem_k_index[231] = 578;
mem_k_index[232] = 581;
mem_k_index[233] = 583;
mem_k_index[234] = 586;
mem_k_index[235] = 588;
mem_k_index[236] = 591;
mem_k_index[237] = 593;
mem_k_index[238] = 596;
mem_k_index[239] = 598;
mem_k_index[240] = 601;
mem_k_index[241] = 603;
mem_k_index[242] = 606;
mem_k_index[243] = 608;
mem_k_index[244] = 611;
mem_k_index[245] = 613;
mem_k_index[246] = 616;
mem_k_index[247] = 618;
mem_k_index[248] = 621;
mem_k_index[249] = 623;
mem_k_index[250] = 626;
mem_k_index[251] = 628;
mem_k_index[252] = 631;
mem_k_index[253] = 633;
mem_k_index[254] = 636;
mem_k_index[255] = 638;
mem_k_index[256] = 960;
mem_k_index[257] = 962;
mem_k_index[258] = 965;
mem_k_index[259] = 967;
mem_k_index[260] = 970;
mem_k_index[261] = 972;
mem_k_index[262] = 975;
mem_k_index[263] = 977;
mem_k_index[264] = 980;
mem_k_index[265] = 982;
mem_k_index[266] = 985;
mem_k_index[267] = 987;
mem_k_index[268] = 990;
mem_k_index[269] = 992;
mem_k_index[270] = 995;
mem_k_index[271] = 997;
mem_k_index[272] = 1000;
mem_k_index[273] = 1002;
mem_k_index[274] = 1005;
mem_k_index[275] = 1007;
mem_k_index[276] = 1010;
mem_k_index[277] = 1012;
mem_k_index[278] = 1015;
mem_k_index[279] = 1017;
mem_k_index[280] = 1020;
mem_k_index[281] = 1022;
mem_k_index[282] = 1025;
mem_k_index[283] = 1027;
mem_k_index[284] = 1030;
mem_k_index[285] = 1032;
mem_k_index[286] = 1035;
mem_k_index[287] = 1037;
mem_k_index[288] = 1040;
mem_k_index[289] = 1042;
mem_k_index[290] = 1045;
mem_k_index[291] = 1047;
mem_k_index[292] = 1050;
mem_k_index[293] = 1052;
mem_k_index[294] = 1055;
mem_k_index[295] = 1057;
mem_k_index[296] = 1060;
mem_k_index[297] = 1062;
mem_k_index[298] = 1065;
mem_k_index[299] = 1068;
mem_k_index[300] = 1070;
mem_k_index[301] = 1073;
mem_k_index[302] = 1075;
mem_k_index[303] = 1078;
mem_k_index[304] = 1080;
mem_k_index[305] = 1083;
mem_k_index[306] = 1085;
mem_k_index[307] = 1088;
mem_k_index[308] = 1090;
mem_k_index[309] = 1093;
mem_k_index[310] = 1095;
mem_k_index[311] = 1098;
mem_k_index[312] = 1100;
mem_k_index[313] = 1103;
mem_k_index[314] = 1105;
mem_k_index[315] = 1108;
mem_k_index[316] = 1110;
mem_k_index[317] = 1113;
mem_k_index[318] = 1115;
mem_k_index[319] = 1118;
mem_k_index[320] = 1120;
mem_k_index[321] = 1123;
mem_k_index[322] = 1125;
mem_k_index[323] = 1128;
mem_k_index[324] = 1130;
mem_k_index[325] = 1133;
mem_k_index[326] = 1135;
mem_k_index[327] = 1138;
mem_k_index[328] = 1140;
mem_k_index[329] = 1143;
mem_k_index[330] = 1145;
mem_k_index[331] = 1148;
mem_k_index[332] = 1150;
mem_k_index[333] = 1153;
mem_k_index[334] = 1155;
mem_k_index[335] = 1158;
mem_k_index[336] = 1160;
mem_k_index[337] = 1163;
mem_k_index[338] = 1165;
mem_k_index[339] = 1168;
mem_k_index[340] = 1170;
mem_k_index[341] = 1173;
mem_k_index[342] = 1176;
mem_k_index[343] = 1178;
mem_k_index[344] = 1181;
mem_k_index[345] = 1183;
mem_k_index[346] = 1186;
mem_k_index[347] = 1188;
mem_k_index[348] = 1191;
mem_k_index[349] = 1193;
mem_k_index[350] = 1196;
mem_k_index[351] = 1198;
mem_k_index[352] = 1201;
mem_k_index[353] = 1203;
mem_k_index[354] = 1206;
mem_k_index[355] = 1208;
mem_k_index[356] = 1211;
mem_k_index[357] = 1213;
mem_k_index[358] = 1216;
mem_k_index[359] = 1218;
mem_k_index[360] = 1221;
mem_k_index[361] = 1223;
mem_k_index[362] = 1226;
mem_k_index[363] = 1228;
mem_k_index[364] = 1231;
mem_k_index[365] = 1233;
mem_k_index[366] = 1236;
mem_k_index[367] = 1238;
mem_k_index[368] = 1241;
mem_k_index[369] = 1243;
mem_k_index[370] = 1246;
mem_k_index[371] = 1248;
mem_k_index[372] = 1251;
mem_k_index[373] = 1253;
mem_k_index[374] = 1256;
mem_k_index[375] = 1258;
mem_k_index[376] = 1261;
mem_k_index[377] = 1263;
mem_k_index[378] = 1266;
mem_k_index[379] = 1268;
mem_k_index[380] = 1271;
mem_k_index[381] = 1273;
mem_k_index[382] = 1276;
mem_k_index[383] = 1278;
mem_k_index[384] = 1600;
mem_k_index[385] = 1602;
mem_k_index[386] = 1605;
mem_k_index[387] = 1607;
mem_k_index[388] = 1610;
mem_k_index[389] = 1612;
mem_k_index[390] = 1615;
mem_k_index[391] = 1617;
mem_k_index[392] = 1620;
mem_k_index[393] = 1622;
mem_k_index[394] = 1625;
mem_k_index[395] = 1627;
mem_k_index[396] = 1630;
mem_k_index[397] = 1632;
mem_k_index[398] = 1635;
mem_k_index[399] = 1637;
mem_k_index[400] = 1640;
mem_k_index[401] = 1642;
mem_k_index[402] = 1645;
mem_k_index[403] = 1647;
mem_k_index[404] = 1650;
mem_k_index[405] = 1652;
mem_k_index[406] = 1655;
mem_k_index[407] = 1657;
mem_k_index[408] = 1660;
mem_k_index[409] = 1662;
mem_k_index[410] = 1665;
mem_k_index[411] = 1667;
mem_k_index[412] = 1670;
mem_k_index[413] = 1672;
mem_k_index[414] = 1675;
mem_k_index[415] = 1677;
mem_k_index[416] = 1680;
mem_k_index[417] = 1682;
mem_k_index[418] = 1685;
mem_k_index[419] = 1687;
mem_k_index[420] = 1690;
mem_k_index[421] = 1692;
mem_k_index[422] = 1695;
mem_k_index[423] = 1697;
mem_k_index[424] = 1700;
mem_k_index[425] = 1702;
mem_k_index[426] = 1705;
mem_k_index[427] = 1708;
mem_k_index[428] = 1710;
mem_k_index[429] = 1713;
mem_k_index[430] = 1715;
mem_k_index[431] = 1718;
mem_k_index[432] = 1720;
mem_k_index[433] = 1723;
mem_k_index[434] = 1725;
mem_k_index[435] = 1728;
mem_k_index[436] = 1730;
mem_k_index[437] = 1733;
mem_k_index[438] = 1735;
mem_k_index[439] = 1738;
mem_k_index[440] = 1740;
mem_k_index[441] = 1743;
mem_k_index[442] = 1745;
mem_k_index[443] = 1748;
mem_k_index[444] = 1750;
mem_k_index[445] = 1753;
mem_k_index[446] = 1755;
mem_k_index[447] = 1758;
mem_k_index[448] = 1760;
mem_k_index[449] = 1763;
mem_k_index[450] = 1765;
mem_k_index[451] = 1768;
mem_k_index[452] = 1770;
mem_k_index[453] = 1773;
mem_k_index[454] = 1775;
mem_k_index[455] = 1778;
mem_k_index[456] = 1780;
mem_k_index[457] = 1783;
mem_k_index[458] = 1785;
mem_k_index[459] = 1788;
mem_k_index[460] = 1790;
mem_k_index[461] = 1793;
mem_k_index[462] = 1795;
mem_k_index[463] = 1798;
mem_k_index[464] = 1800;
mem_k_index[465] = 1803;
mem_k_index[466] = 1805;
mem_k_index[467] = 1808;
mem_k_index[468] = 1810;
mem_k_index[469] = 1813;
mem_k_index[470] = 1816;
mem_k_index[471] = 1818;
mem_k_index[472] = 1821;
mem_k_index[473] = 1823;
mem_k_index[474] = 1826;
mem_k_index[475] = 1828;
mem_k_index[476] = 1831;
mem_k_index[477] = 1833;
mem_k_index[478] = 1836;
mem_k_index[479] = 1838;
mem_k_index[480] = 1841;
mem_k_index[481] = 1843;
mem_k_index[482] = 1846;
mem_k_index[483] = 1848;
mem_k_index[484] = 1851;
mem_k_index[485] = 1853;
mem_k_index[486] = 1856;
mem_k_index[487] = 1858;
mem_k_index[488] = 1861;
mem_k_index[489] = 1863;
mem_k_index[490] = 1866;
mem_k_index[491] = 1868;
mem_k_index[492] = 1871;
mem_k_index[493] = 1873;
mem_k_index[494] = 1876;
mem_k_index[495] = 1878;
mem_k_index[496] = 1881;
mem_k_index[497] = 1883;
mem_k_index[498] = 1886;
mem_k_index[499] = 1888;
mem_k_index[500] = 1891;
mem_k_index[501] = 1893;
mem_k_index[502] = 1896;
mem_k_index[503] = 1898;
mem_k_index[504] = 1901;
mem_k_index[505] = 1903;
mem_k_index[506] = 1906;
mem_k_index[507] = 1908;
mem_k_index[508] = 1911;
mem_k_index[509] = 1913;
mem_k_index[510] = 1916;
mem_k_index[511] = 1918;
mem_k_index[512] = 2240;
mem_k_index[513] = 2242;
mem_k_index[514] = 2245;
mem_k_index[515] = 2247;
mem_k_index[516] = 2250;
mem_k_index[517] = 2252;
mem_k_index[518] = 2255;
mem_k_index[519] = 2257;
mem_k_index[520] = 2260;
mem_k_index[521] = 2262;
mem_k_index[522] = 2265;
mem_k_index[523] = 2267;
mem_k_index[524] = 2270;
mem_k_index[525] = 2272;
mem_k_index[526] = 2275;
mem_k_index[527] = 2277;
mem_k_index[528] = 2280;
mem_k_index[529] = 2282;
mem_k_index[530] = 2285;
mem_k_index[531] = 2287;
mem_k_index[532] = 2290;
mem_k_index[533] = 2292;
mem_k_index[534] = 2295;
mem_k_index[535] = 2297;
mem_k_index[536] = 2300;
mem_k_index[537] = 2302;
mem_k_index[538] = 2305;
mem_k_index[539] = 2307;
mem_k_index[540] = 2310;
mem_k_index[541] = 2312;
mem_k_index[542] = 2315;
mem_k_index[543] = 2317;
mem_k_index[544] = 2320;
mem_k_index[545] = 2322;
mem_k_index[546] = 2325;
mem_k_index[547] = 2327;
mem_k_index[548] = 2330;
mem_k_index[549] = 2332;
mem_k_index[550] = 2335;
mem_k_index[551] = 2337;
mem_k_index[552] = 2340;
mem_k_index[553] = 2342;
mem_k_index[554] = 2345;
mem_k_index[555] = 2348;
mem_k_index[556] = 2350;
mem_k_index[557] = 2353;
mem_k_index[558] = 2355;
mem_k_index[559] = 2358;
mem_k_index[560] = 2360;
mem_k_index[561] = 2363;
mem_k_index[562] = 2365;
mem_k_index[563] = 2368;
mem_k_index[564] = 2370;
mem_k_index[565] = 2373;
mem_k_index[566] = 2375;
mem_k_index[567] = 2378;
mem_k_index[568] = 2380;
mem_k_index[569] = 2383;
mem_k_index[570] = 2385;
mem_k_index[571] = 2388;
mem_k_index[572] = 2390;
mem_k_index[573] = 2393;
mem_k_index[574] = 2395;
mem_k_index[575] = 2398;
mem_k_index[576] = 2400;
mem_k_index[577] = 2403;
mem_k_index[578] = 2405;
mem_k_index[579] = 2408;
mem_k_index[580] = 2410;
mem_k_index[581] = 2413;
mem_k_index[582] = 2415;
mem_k_index[583] = 2418;
mem_k_index[584] = 2420;
mem_k_index[585] = 2423;
mem_k_index[586] = 2425;
mem_k_index[587] = 2428;
mem_k_index[588] = 2430;
mem_k_index[589] = 2433;
mem_k_index[590] = 2435;
mem_k_index[591] = 2438;
mem_k_index[592] = 2440;
mem_k_index[593] = 2443;
mem_k_index[594] = 2445;
mem_k_index[595] = 2448;
mem_k_index[596] = 2450;
mem_k_index[597] = 2453;
mem_k_index[598] = 2456;
mem_k_index[599] = 2458;
mem_k_index[600] = 2461;
mem_k_index[601] = 2463;
mem_k_index[602] = 2466;
mem_k_index[603] = 2468;
mem_k_index[604] = 2471;
mem_k_index[605] = 2473;
mem_k_index[606] = 2476;
mem_k_index[607] = 2478;
mem_k_index[608] = 2481;
mem_k_index[609] = 2483;
mem_k_index[610] = 2486;
mem_k_index[611] = 2488;
mem_k_index[612] = 2491;
mem_k_index[613] = 2493;
mem_k_index[614] = 2496;
mem_k_index[615] = 2498;
mem_k_index[616] = 2501;
mem_k_index[617] = 2503;
mem_k_index[618] = 2506;
mem_k_index[619] = 2508;
mem_k_index[620] = 2511;
mem_k_index[621] = 2513;
mem_k_index[622] = 2516;
mem_k_index[623] = 2518;
mem_k_index[624] = 2521;
mem_k_index[625] = 2523;
mem_k_index[626] = 2526;
mem_k_index[627] = 2528;
mem_k_index[628] = 2531;
mem_k_index[629] = 2533;
mem_k_index[630] = 2536;
mem_k_index[631] = 2538;
mem_k_index[632] = 2541;
mem_k_index[633] = 2543;
mem_k_index[634] = 2546;
mem_k_index[635] = 2548;
mem_k_index[636] = 2551;
mem_k_index[637] = 2553;
mem_k_index[638] = 2556;
mem_k_index[639] = 2558;
mem_k_index[640] = 2880;
mem_k_index[641] = 2882;
mem_k_index[642] = 2885;
mem_k_index[643] = 2887;
mem_k_index[644] = 2890;
mem_k_index[645] = 2892;
mem_k_index[646] = 2895;
mem_k_index[647] = 2897;
mem_k_index[648] = 2900;
mem_k_index[649] = 2902;
mem_k_index[650] = 2905;
mem_k_index[651] = 2907;
mem_k_index[652] = 2910;
mem_k_index[653] = 2912;
mem_k_index[654] = 2915;
mem_k_index[655] = 2917;
mem_k_index[656] = 2920;
mem_k_index[657] = 2922;
mem_k_index[658] = 2925;
mem_k_index[659] = 2927;
mem_k_index[660] = 2930;
mem_k_index[661] = 2932;
mem_k_index[662] = 2935;
mem_k_index[663] = 2937;
mem_k_index[664] = 2940;
mem_k_index[665] = 2942;
mem_k_index[666] = 2945;
mem_k_index[667] = 2947;
mem_k_index[668] = 2950;
mem_k_index[669] = 2952;
mem_k_index[670] = 2955;
mem_k_index[671] = 2957;
mem_k_index[672] = 2960;
mem_k_index[673] = 2962;
mem_k_index[674] = 2965;
mem_k_index[675] = 2967;
mem_k_index[676] = 2970;
mem_k_index[677] = 2972;
mem_k_index[678] = 2975;
mem_k_index[679] = 2977;
mem_k_index[680] = 2980;
mem_k_index[681] = 2982;
mem_k_index[682] = 2985;
mem_k_index[683] = 2988;
mem_k_index[684] = 2990;
mem_k_index[685] = 2993;
mem_k_index[686] = 2995;
mem_k_index[687] = 2998;
mem_k_index[688] = 3000;
mem_k_index[689] = 3003;
mem_k_index[690] = 3005;
mem_k_index[691] = 3008;
mem_k_index[692] = 3010;
mem_k_index[693] = 3013;
mem_k_index[694] = 3015;
mem_k_index[695] = 3018;
mem_k_index[696] = 3020;
mem_k_index[697] = 3023;
mem_k_index[698] = 3025;
mem_k_index[699] = 3028;
mem_k_index[700] = 3030;
mem_k_index[701] = 3033;
mem_k_index[702] = 3035;
mem_k_index[703] = 3038;
mem_k_index[704] = 3040;
mem_k_index[705] = 3043;
mem_k_index[706] = 3045;
mem_k_index[707] = 3048;
mem_k_index[708] = 3050;
mem_k_index[709] = 3053;
mem_k_index[710] = 3055;
mem_k_index[711] = 3058;
mem_k_index[712] = 3060;
mem_k_index[713] = 3063;
mem_k_index[714] = 3065;
mem_k_index[715] = 3068;
mem_k_index[716] = 3070;
mem_k_index[717] = 3073;
mem_k_index[718] = 3075;
mem_k_index[719] = 3078;
mem_k_index[720] = 3080;
mem_k_index[721] = 3083;
mem_k_index[722] = 3085;
mem_k_index[723] = 3088;
mem_k_index[724] = 3090;
mem_k_index[725] = 3093;
mem_k_index[726] = 3096;
mem_k_index[727] = 3098;
mem_k_index[728] = 3101;
mem_k_index[729] = 3103;
mem_k_index[730] = 3106;
mem_k_index[731] = 3108;
mem_k_index[732] = 3111;
mem_k_index[733] = 3113;
mem_k_index[734] = 3116;
mem_k_index[735] = 3118;
mem_k_index[736] = 3121;
mem_k_index[737] = 3123;
mem_k_index[738] = 3126;
mem_k_index[739] = 3128;
mem_k_index[740] = 3131;
mem_k_index[741] = 3133;
mem_k_index[742] = 3136;
mem_k_index[743] = 3138;
mem_k_index[744] = 3141;
mem_k_index[745] = 3143;
mem_k_index[746] = 3146;
mem_k_index[747] = 3148;
mem_k_index[748] = 3151;
mem_k_index[749] = 3153;
mem_k_index[750] = 3156;
mem_k_index[751] = 3158;
mem_k_index[752] = 3161;
mem_k_index[753] = 3163;
mem_k_index[754] = 3166;
mem_k_index[755] = 3168;
mem_k_index[756] = 3171;
mem_k_index[757] = 3173;
mem_k_index[758] = 3176;
mem_k_index[759] = 3178;
mem_k_index[760] = 3181;
mem_k_index[761] = 3183;
mem_k_index[762] = 3186;
mem_k_index[763] = 3188;
mem_k_index[764] = 3191;
mem_k_index[765] = 3193;
mem_k_index[766] = 3196;
mem_k_index[767] = 3198;
mem_k_index[768] = 3520;
mem_k_index[769] = 3522;
mem_k_index[770] = 3525;
mem_k_index[771] = 3527;
mem_k_index[772] = 3530;
mem_k_index[773] = 3532;
mem_k_index[774] = 3535;
mem_k_index[775] = 3537;
mem_k_index[776] = 3540;
mem_k_index[777] = 3542;
mem_k_index[778] = 3545;
mem_k_index[779] = 3547;
mem_k_index[780] = 3550;
mem_k_index[781] = 3552;
mem_k_index[782] = 3555;
mem_k_index[783] = 3557;
mem_k_index[784] = 3560;
mem_k_index[785] = 3562;
mem_k_index[786] = 3565;
mem_k_index[787] = 3567;
mem_k_index[788] = 3570;
mem_k_index[789] = 3572;
mem_k_index[790] = 3575;
mem_k_index[791] = 3577;
mem_k_index[792] = 3580;
mem_k_index[793] = 3582;
mem_k_index[794] = 3585;
mem_k_index[795] = 3587;
mem_k_index[796] = 3590;
mem_k_index[797] = 3592;
mem_k_index[798] = 3595;
mem_k_index[799] = 3597;
mem_k_index[800] = 3600;
mem_k_index[801] = 3602;
mem_k_index[802] = 3605;
mem_k_index[803] = 3607;
mem_k_index[804] = 3610;
mem_k_index[805] = 3612;
mem_k_index[806] = 3615;
mem_k_index[807] = 3617;
mem_k_index[808] = 3620;
mem_k_index[809] = 3622;
mem_k_index[810] = 3625;
mem_k_index[811] = 3628;
mem_k_index[812] = 3630;
mem_k_index[813] = 3633;
mem_k_index[814] = 3635;
mem_k_index[815] = 3638;
mem_k_index[816] = 3640;
mem_k_index[817] = 3643;
mem_k_index[818] = 3645;
mem_k_index[819] = 3648;
mem_k_index[820] = 3650;
mem_k_index[821] = 3653;
mem_k_index[822] = 3655;
mem_k_index[823] = 3658;
mem_k_index[824] = 3660;
mem_k_index[825] = 3663;
mem_k_index[826] = 3665;
mem_k_index[827] = 3668;
mem_k_index[828] = 3670;
mem_k_index[829] = 3673;
mem_k_index[830] = 3675;
mem_k_index[831] = 3678;
mem_k_index[832] = 3680;
mem_k_index[833] = 3683;
mem_k_index[834] = 3685;
mem_k_index[835] = 3688;
mem_k_index[836] = 3690;
mem_k_index[837] = 3693;
mem_k_index[838] = 3695;
mem_k_index[839] = 3698;
mem_k_index[840] = 3700;
mem_k_index[841] = 3703;
mem_k_index[842] = 3705;
mem_k_index[843] = 3708;
mem_k_index[844] = 3710;
mem_k_index[845] = 3713;
mem_k_index[846] = 3715;
mem_k_index[847] = 3718;
mem_k_index[848] = 3720;
mem_k_index[849] = 3723;
mem_k_index[850] = 3725;
mem_k_index[851] = 3728;
mem_k_index[852] = 3730;
mem_k_index[853] = 3733;
mem_k_index[854] = 3736;
mem_k_index[855] = 3738;
mem_k_index[856] = 3741;
mem_k_index[857] = 3743;
mem_k_index[858] = 3746;
mem_k_index[859] = 3748;
mem_k_index[860] = 3751;
mem_k_index[861] = 3753;
mem_k_index[862] = 3756;
mem_k_index[863] = 3758;
mem_k_index[864] = 3761;
mem_k_index[865] = 3763;
mem_k_index[866] = 3766;
mem_k_index[867] = 3768;
mem_k_index[868] = 3771;
mem_k_index[869] = 3773;
mem_k_index[870] = 3776;
mem_k_index[871] = 3778;
mem_k_index[872] = 3781;
mem_k_index[873] = 3783;
mem_k_index[874] = 3786;
mem_k_index[875] = 3788;
mem_k_index[876] = 3791;
mem_k_index[877] = 3793;
mem_k_index[878] = 3796;
mem_k_index[879] = 3798;
mem_k_index[880] = 3801;
mem_k_index[881] = 3803;
mem_k_index[882] = 3806;
mem_k_index[883] = 3808;
mem_k_index[884] = 3811;
mem_k_index[885] = 3813;
mem_k_index[886] = 3816;
mem_k_index[887] = 3818;
mem_k_index[888] = 3821;
mem_k_index[889] = 3823;
mem_k_index[890] = 3826;
mem_k_index[891] = 3828;
mem_k_index[892] = 3831;
mem_k_index[893] = 3833;
mem_k_index[894] = 3836;
mem_k_index[895] = 3838;
mem_k_index[896] = 4160;
mem_k_index[897] = 4162;
mem_k_index[898] = 4165;
mem_k_index[899] = 4167;
mem_k_index[900] = 4170;
mem_k_index[901] = 4172;
mem_k_index[902] = 4175;
mem_k_index[903] = 4177;
mem_k_index[904] = 4180;
mem_k_index[905] = 4182;
mem_k_index[906] = 4185;
mem_k_index[907] = 4187;
mem_k_index[908] = 4190;
mem_k_index[909] = 4192;
mem_k_index[910] = 4195;
mem_k_index[911] = 4197;
mem_k_index[912] = 4200;
mem_k_index[913] = 4202;
mem_k_index[914] = 4205;
mem_k_index[915] = 4207;
mem_k_index[916] = 4210;
mem_k_index[917] = 4212;
mem_k_index[918] = 4215;
mem_k_index[919] = 4217;
mem_k_index[920] = 4220;
mem_k_index[921] = 4222;
mem_k_index[922] = 4225;
mem_k_index[923] = 4227;
mem_k_index[924] = 4230;
mem_k_index[925] = 4232;
mem_k_index[926] = 4235;
mem_k_index[927] = 4237;
mem_k_index[928] = 4240;
mem_k_index[929] = 4242;
mem_k_index[930] = 4245;
mem_k_index[931] = 4247;
mem_k_index[932] = 4250;
mem_k_index[933] = 4252;
mem_k_index[934] = 4255;
mem_k_index[935] = 4257;
mem_k_index[936] = 4260;
mem_k_index[937] = 4262;
mem_k_index[938] = 4265;
mem_k_index[939] = 4268;
mem_k_index[940] = 4270;
mem_k_index[941] = 4273;
mem_k_index[942] = 4275;
mem_k_index[943] = 4278;
mem_k_index[944] = 4280;
mem_k_index[945] = 4283;
mem_k_index[946] = 4285;
mem_k_index[947] = 4288;
mem_k_index[948] = 4290;
mem_k_index[949] = 4293;
mem_k_index[950] = 4295;
mem_k_index[951] = 4298;
mem_k_index[952] = 4300;
mem_k_index[953] = 4303;
mem_k_index[954] = 4305;
mem_k_index[955] = 4308;
mem_k_index[956] = 4310;
mem_k_index[957] = 4313;
mem_k_index[958] = 4315;
mem_k_index[959] = 4318;
mem_k_index[960] = 4320;
mem_k_index[961] = 4323;
mem_k_index[962] = 4325;
mem_k_index[963] = 4328;
mem_k_index[964] = 4330;
mem_k_index[965] = 4333;
mem_k_index[966] = 4335;
mem_k_index[967] = 4338;
mem_k_index[968] = 4340;
mem_k_index[969] = 4343;
mem_k_index[970] = 4345;
mem_k_index[971] = 4348;
mem_k_index[972] = 4350;
mem_k_index[973] = 4353;
mem_k_index[974] = 4355;
mem_k_index[975] = 4358;
mem_k_index[976] = 4360;
mem_k_index[977] = 4363;
mem_k_index[978] = 4365;
mem_k_index[979] = 4368;
mem_k_index[980] = 4370;
mem_k_index[981] = 4373;
mem_k_index[982] = 4376;
mem_k_index[983] = 4378;
mem_k_index[984] = 4381;
mem_k_index[985] = 4383;
mem_k_index[986] = 4386;
mem_k_index[987] = 4388;
mem_k_index[988] = 4391;
mem_k_index[989] = 4393;
mem_k_index[990] = 4396;
mem_k_index[991] = 4398;
mem_k_index[992] = 4401;
mem_k_index[993] = 4403;
mem_k_index[994] = 4406;
mem_k_index[995] = 4408;
mem_k_index[996] = 4411;
mem_k_index[997] = 4413;
mem_k_index[998] = 4416;
mem_k_index[999] = 4418;
mem_k_index[1000] = 4421;
mem_k_index[1001] = 4423;
mem_k_index[1002] = 4426;
mem_k_index[1003] = 4428;
mem_k_index[1004] = 4431;
mem_k_index[1005] = 4433;
mem_k_index[1006] = 4436;
mem_k_index[1007] = 4438;
mem_k_index[1008] = 4441;
mem_k_index[1009] = 4443;
mem_k_index[1010] = 4446;
mem_k_index[1011] = 4448;
mem_k_index[1012] = 4451;
mem_k_index[1013] = 4453;
mem_k_index[1014] = 4456;
mem_k_index[1015] = 4458;
mem_k_index[1016] = 4461;
mem_k_index[1017] = 4463;
mem_k_index[1018] = 4466;
mem_k_index[1019] = 4468;
mem_k_index[1020] = 4471;
mem_k_index[1021] = 4473;
mem_k_index[1022] = 4476;
mem_k_index[1023] = 4478;
mem_k_index[1024] = 4800;
mem_k_index[1025] = 4802;
mem_k_index[1026] = 4805;
mem_k_index[1027] = 4807;
mem_k_index[1028] = 4810;
mem_k_index[1029] = 4812;
mem_k_index[1030] = 4815;
mem_k_index[1031] = 4817;
mem_k_index[1032] = 4820;
mem_k_index[1033] = 4822;
mem_k_index[1034] = 4825;
mem_k_index[1035] = 4827;
mem_k_index[1036] = 4830;
mem_k_index[1037] = 4832;
mem_k_index[1038] = 4835;
mem_k_index[1039] = 4837;
mem_k_index[1040] = 4840;
mem_k_index[1041] = 4842;
mem_k_index[1042] = 4845;
mem_k_index[1043] = 4847;
mem_k_index[1044] = 4850;
mem_k_index[1045] = 4852;
mem_k_index[1046] = 4855;
mem_k_index[1047] = 4857;
mem_k_index[1048] = 4860;
mem_k_index[1049] = 4862;
mem_k_index[1050] = 4865;
mem_k_index[1051] = 4867;
mem_k_index[1052] = 4870;
mem_k_index[1053] = 4872;
mem_k_index[1054] = 4875;
mem_k_index[1055] = 4877;
mem_k_index[1056] = 4880;
mem_k_index[1057] = 4882;
mem_k_index[1058] = 4885;
mem_k_index[1059] = 4887;
mem_k_index[1060] = 4890;
mem_k_index[1061] = 4892;
mem_k_index[1062] = 4895;
mem_k_index[1063] = 4897;
mem_k_index[1064] = 4900;
mem_k_index[1065] = 4902;
mem_k_index[1066] = 4905;
mem_k_index[1067] = 4908;
mem_k_index[1068] = 4910;
mem_k_index[1069] = 4913;
mem_k_index[1070] = 4915;
mem_k_index[1071] = 4918;
mem_k_index[1072] = 4920;
mem_k_index[1073] = 4923;
mem_k_index[1074] = 4925;
mem_k_index[1075] = 4928;
mem_k_index[1076] = 4930;
mem_k_index[1077] = 4933;
mem_k_index[1078] = 4935;
mem_k_index[1079] = 4938;
mem_k_index[1080] = 4940;
mem_k_index[1081] = 4943;
mem_k_index[1082] = 4945;
mem_k_index[1083] = 4948;
mem_k_index[1084] = 4950;
mem_k_index[1085] = 4953;
mem_k_index[1086] = 4955;
mem_k_index[1087] = 4958;
mem_k_index[1088] = 4960;
mem_k_index[1089] = 4963;
mem_k_index[1090] = 4965;
mem_k_index[1091] = 4968;
mem_k_index[1092] = 4970;
mem_k_index[1093] = 4973;
mem_k_index[1094] = 4975;
mem_k_index[1095] = 4978;
mem_k_index[1096] = 4980;
mem_k_index[1097] = 4983;
mem_k_index[1098] = 4985;
mem_k_index[1099] = 4988;
mem_k_index[1100] = 4990;
mem_k_index[1101] = 4993;
mem_k_index[1102] = 4995;
mem_k_index[1103] = 4998;
mem_k_index[1104] = 5000;
mem_k_index[1105] = 5003;
mem_k_index[1106] = 5005;
mem_k_index[1107] = 5008;
mem_k_index[1108] = 5010;
mem_k_index[1109] = 5013;
mem_k_index[1110] = 5016;
mem_k_index[1111] = 5018;
mem_k_index[1112] = 5021;
mem_k_index[1113] = 5023;
mem_k_index[1114] = 5026;
mem_k_index[1115] = 5028;
mem_k_index[1116] = 5031;
mem_k_index[1117] = 5033;
mem_k_index[1118] = 5036;
mem_k_index[1119] = 5038;
mem_k_index[1120] = 5041;
mem_k_index[1121] = 5043;
mem_k_index[1122] = 5046;
mem_k_index[1123] = 5048;
mem_k_index[1124] = 5051;
mem_k_index[1125] = 5053;
mem_k_index[1126] = 5056;
mem_k_index[1127] = 5058;
mem_k_index[1128] = 5061;
mem_k_index[1129] = 5063;
mem_k_index[1130] = 5066;
mem_k_index[1131] = 5068;
mem_k_index[1132] = 5071;
mem_k_index[1133] = 5073;
mem_k_index[1134] = 5076;
mem_k_index[1135] = 5078;
mem_k_index[1136] = 5081;
mem_k_index[1137] = 5083;
mem_k_index[1138] = 5086;
mem_k_index[1139] = 5088;
mem_k_index[1140] = 5091;
mem_k_index[1141] = 5093;
mem_k_index[1142] = 5096;
mem_k_index[1143] = 5098;
mem_k_index[1144] = 5101;
mem_k_index[1145] = 5103;
mem_k_index[1146] = 5106;
mem_k_index[1147] = 5108;
mem_k_index[1148] = 5111;
mem_k_index[1149] = 5113;
mem_k_index[1150] = 5116;
mem_k_index[1151] = 5118;
mem_k_index[1152] = 5120;
mem_k_index[1153] = 5122;
mem_k_index[1154] = 5125;
mem_k_index[1155] = 5127;
mem_k_index[1156] = 5130;
mem_k_index[1157] = 5132;
mem_k_index[1158] = 5135;
mem_k_index[1159] = 5137;
mem_k_index[1160] = 5140;
mem_k_index[1161] = 5142;
mem_k_index[1162] = 5145;
mem_k_index[1163] = 5147;
mem_k_index[1164] = 5150;
mem_k_index[1165] = 5152;
mem_k_index[1166] = 5155;
mem_k_index[1167] = 5157;
mem_k_index[1168] = 5160;
mem_k_index[1169] = 5162;
mem_k_index[1170] = 5165;
mem_k_index[1171] = 5167;
mem_k_index[1172] = 5170;
mem_k_index[1173] = 5172;
mem_k_index[1174] = 5175;
mem_k_index[1175] = 5177;
mem_k_index[1176] = 5180;
mem_k_index[1177] = 5182;
mem_k_index[1178] = 5185;
mem_k_index[1179] = 5187;
mem_k_index[1180] = 5190;
mem_k_index[1181] = 5192;
mem_k_index[1182] = 5195;
mem_k_index[1183] = 5197;
mem_k_index[1184] = 5200;
mem_k_index[1185] = 5202;
mem_k_index[1186] = 5205;
mem_k_index[1187] = 5207;
mem_k_index[1188] = 5210;
mem_k_index[1189] = 5212;
mem_k_index[1190] = 5215;
mem_k_index[1191] = 5217;
mem_k_index[1192] = 5220;
mem_k_index[1193] = 5222;
mem_k_index[1194] = 5225;
mem_k_index[1195] = 5228;
mem_k_index[1196] = 5230;
mem_k_index[1197] = 5233;
mem_k_index[1198] = 5235;
mem_k_index[1199] = 5238;
mem_k_index[1200] = 5240;
mem_k_index[1201] = 5243;
mem_k_index[1202] = 5245;
mem_k_index[1203] = 5248;
mem_k_index[1204] = 5250;
mem_k_index[1205] = 5253;
mem_k_index[1206] = 5255;
mem_k_index[1207] = 5258;
mem_k_index[1208] = 5260;
mem_k_index[1209] = 5263;
mem_k_index[1210] = 5265;
mem_k_index[1211] = 5268;
mem_k_index[1212] = 5270;
mem_k_index[1213] = 5273;
mem_k_index[1214] = 5275;
mem_k_index[1215] = 5278;
mem_k_index[1216] = 5280;
mem_k_index[1217] = 5283;
mem_k_index[1218] = 5285;
mem_k_index[1219] = 5288;
mem_k_index[1220] = 5290;
mem_k_index[1221] = 5293;
mem_k_index[1222] = 5295;
mem_k_index[1223] = 5298;
mem_k_index[1224] = 5300;
mem_k_index[1225] = 5303;
mem_k_index[1226] = 5305;
mem_k_index[1227] = 5308;
mem_k_index[1228] = 5310;
mem_k_index[1229] = 5313;
mem_k_index[1230] = 5315;
mem_k_index[1231] = 5318;
mem_k_index[1232] = 5320;
mem_k_index[1233] = 5323;
mem_k_index[1234] = 5325;
mem_k_index[1235] = 5328;
mem_k_index[1236] = 5330;
mem_k_index[1237] = 5333;
mem_k_index[1238] = 5336;
mem_k_index[1239] = 5338;
mem_k_index[1240] = 5341;
mem_k_index[1241] = 5343;
mem_k_index[1242] = 5346;
mem_k_index[1243] = 5348;
mem_k_index[1244] = 5351;
mem_k_index[1245] = 5353;
mem_k_index[1246] = 5356;
mem_k_index[1247] = 5358;
mem_k_index[1248] = 5361;
mem_k_index[1249] = 5363;
mem_k_index[1250] = 5366;
mem_k_index[1251] = 5368;
mem_k_index[1252] = 5371;
mem_k_index[1253] = 5373;
mem_k_index[1254] = 5376;
mem_k_index[1255] = 5378;
mem_k_index[1256] = 5381;
mem_k_index[1257] = 5383;
mem_k_index[1258] = 5386;
mem_k_index[1259] = 5388;
mem_k_index[1260] = 5391;
mem_k_index[1261] = 5393;
mem_k_index[1262] = 5396;
mem_k_index[1263] = 5398;
mem_k_index[1264] = 5401;
mem_k_index[1265] = 5403;
mem_k_index[1266] = 5406;
mem_k_index[1267] = 5408;
mem_k_index[1268] = 5411;
mem_k_index[1269] = 5413;
mem_k_index[1270] = 5416;
mem_k_index[1271] = 5418;
mem_k_index[1272] = 5421;
mem_k_index[1273] = 5423;
mem_k_index[1274] = 5426;
mem_k_index[1275] = 5428;
mem_k_index[1276] = 5431;
mem_k_index[1277] = 5433;
mem_k_index[1278] = 5436;
mem_k_index[1279] = 5438;
mem_k_index[1280] = 5760;
mem_k_index[1281] = 5762;
mem_k_index[1282] = 5765;
mem_k_index[1283] = 5767;
mem_k_index[1284] = 5770;
mem_k_index[1285] = 5772;
mem_k_index[1286] = 5775;
mem_k_index[1287] = 5777;
mem_k_index[1288] = 5780;
mem_k_index[1289] = 5782;
mem_k_index[1290] = 5785;
mem_k_index[1291] = 5787;
mem_k_index[1292] = 5790;
mem_k_index[1293] = 5792;
mem_k_index[1294] = 5795;
mem_k_index[1295] = 5797;
mem_k_index[1296] = 5800;
mem_k_index[1297] = 5802;
mem_k_index[1298] = 5805;
mem_k_index[1299] = 5807;
mem_k_index[1300] = 5810;
mem_k_index[1301] = 5812;
mem_k_index[1302] = 5815;
mem_k_index[1303] = 5817;
mem_k_index[1304] = 5820;
mem_k_index[1305] = 5822;
mem_k_index[1306] = 5825;
mem_k_index[1307] = 5827;
mem_k_index[1308] = 5830;
mem_k_index[1309] = 5832;
mem_k_index[1310] = 5835;
mem_k_index[1311] = 5837;
mem_k_index[1312] = 5840;
mem_k_index[1313] = 5842;
mem_k_index[1314] = 5845;
mem_k_index[1315] = 5847;
mem_k_index[1316] = 5850;
mem_k_index[1317] = 5852;
mem_k_index[1318] = 5855;
mem_k_index[1319] = 5857;
mem_k_index[1320] = 5860;
mem_k_index[1321] = 5862;
mem_k_index[1322] = 5865;
mem_k_index[1323] = 5868;
mem_k_index[1324] = 5870;
mem_k_index[1325] = 5873;
mem_k_index[1326] = 5875;
mem_k_index[1327] = 5878;
mem_k_index[1328] = 5880;
mem_k_index[1329] = 5883;
mem_k_index[1330] = 5885;
mem_k_index[1331] = 5888;
mem_k_index[1332] = 5890;
mem_k_index[1333] = 5893;
mem_k_index[1334] = 5895;
mem_k_index[1335] = 5898;
mem_k_index[1336] = 5900;
mem_k_index[1337] = 5903;
mem_k_index[1338] = 5905;
mem_k_index[1339] = 5908;
mem_k_index[1340] = 5910;
mem_k_index[1341] = 5913;
mem_k_index[1342] = 5915;
mem_k_index[1343] = 5918;
mem_k_index[1344] = 5920;
mem_k_index[1345] = 5923;
mem_k_index[1346] = 5925;
mem_k_index[1347] = 5928;
mem_k_index[1348] = 5930;
mem_k_index[1349] = 5933;
mem_k_index[1350] = 5935;
mem_k_index[1351] = 5938;
mem_k_index[1352] = 5940;
mem_k_index[1353] = 5943;
mem_k_index[1354] = 5945;
mem_k_index[1355] = 5948;
mem_k_index[1356] = 5950;
mem_k_index[1357] = 5953;
mem_k_index[1358] = 5955;
mem_k_index[1359] = 5958;
mem_k_index[1360] = 5960;
mem_k_index[1361] = 5963;
mem_k_index[1362] = 5965;
mem_k_index[1363] = 5968;
mem_k_index[1364] = 5970;
mem_k_index[1365] = 5973;
mem_k_index[1366] = 5976;
mem_k_index[1367] = 5978;
mem_k_index[1368] = 5981;
mem_k_index[1369] = 5983;
mem_k_index[1370] = 5986;
mem_k_index[1371] = 5988;
mem_k_index[1372] = 5991;
mem_k_index[1373] = 5993;
mem_k_index[1374] = 5996;
mem_k_index[1375] = 5998;
mem_k_index[1376] = 6001;
mem_k_index[1377] = 6003;
mem_k_index[1378] = 6006;
mem_k_index[1379] = 6008;
mem_k_index[1380] = 6011;
mem_k_index[1381] = 6013;
mem_k_index[1382] = 6016;
mem_k_index[1383] = 6018;
mem_k_index[1384] = 6021;
mem_k_index[1385] = 6023;
mem_k_index[1386] = 6026;
mem_k_index[1387] = 6028;
mem_k_index[1388] = 6031;
mem_k_index[1389] = 6033;
mem_k_index[1390] = 6036;
mem_k_index[1391] = 6038;
mem_k_index[1392] = 6041;
mem_k_index[1393] = 6043;
mem_k_index[1394] = 6046;
mem_k_index[1395] = 6048;
mem_k_index[1396] = 6051;
mem_k_index[1397] = 6053;
mem_k_index[1398] = 6056;
mem_k_index[1399] = 6058;
mem_k_index[1400] = 6061;
mem_k_index[1401] = 6063;
mem_k_index[1402] = 6066;
mem_k_index[1403] = 6068;
mem_k_index[1404] = 6071;
mem_k_index[1405] = 6073;
mem_k_index[1406] = 6076;
mem_k_index[1407] = 6078;
mem_k_index[1408] = 6400;
mem_k_index[1409] = 6402;
mem_k_index[1410] = 6405;
mem_k_index[1411] = 6407;
mem_k_index[1412] = 6410;
mem_k_index[1413] = 6412;
mem_k_index[1414] = 6415;
mem_k_index[1415] = 6417;
mem_k_index[1416] = 6420;
mem_k_index[1417] = 6422;
mem_k_index[1418] = 6425;
mem_k_index[1419] = 6427;
mem_k_index[1420] = 6430;
mem_k_index[1421] = 6432;
mem_k_index[1422] = 6435;
mem_k_index[1423] = 6437;
mem_k_index[1424] = 6440;
mem_k_index[1425] = 6442;
mem_k_index[1426] = 6445;
mem_k_index[1427] = 6447;
mem_k_index[1428] = 6450;
mem_k_index[1429] = 6452;
mem_k_index[1430] = 6455;
mem_k_index[1431] = 6457;
mem_k_index[1432] = 6460;
mem_k_index[1433] = 6462;
mem_k_index[1434] = 6465;
mem_k_index[1435] = 6467;
mem_k_index[1436] = 6470;
mem_k_index[1437] = 6472;
mem_k_index[1438] = 6475;
mem_k_index[1439] = 6477;
mem_k_index[1440] = 6480;
mem_k_index[1441] = 6482;
mem_k_index[1442] = 6485;
mem_k_index[1443] = 6487;
mem_k_index[1444] = 6490;
mem_k_index[1445] = 6492;
mem_k_index[1446] = 6495;
mem_k_index[1447] = 6497;
mem_k_index[1448] = 6500;
mem_k_index[1449] = 6502;
mem_k_index[1450] = 6505;
mem_k_index[1451] = 6508;
mem_k_index[1452] = 6510;
mem_k_index[1453] = 6513;
mem_k_index[1454] = 6515;
mem_k_index[1455] = 6518;
mem_k_index[1456] = 6520;
mem_k_index[1457] = 6523;
mem_k_index[1458] = 6525;
mem_k_index[1459] = 6528;
mem_k_index[1460] = 6530;
mem_k_index[1461] = 6533;
mem_k_index[1462] = 6535;
mem_k_index[1463] = 6538;
mem_k_index[1464] = 6540;
mem_k_index[1465] = 6543;
mem_k_index[1466] = 6545;
mem_k_index[1467] = 6548;
mem_k_index[1468] = 6550;
mem_k_index[1469] = 6553;
mem_k_index[1470] = 6555;
mem_k_index[1471] = 6558;
mem_k_index[1472] = 6560;
mem_k_index[1473] = 6563;
mem_k_index[1474] = 6565;
mem_k_index[1475] = 6568;
mem_k_index[1476] = 6570;
mem_k_index[1477] = 6573;
mem_k_index[1478] = 6575;
mem_k_index[1479] = 6578;
mem_k_index[1480] = 6580;
mem_k_index[1481] = 6583;
mem_k_index[1482] = 6585;
mem_k_index[1483] = 6588;
mem_k_index[1484] = 6590;
mem_k_index[1485] = 6593;
mem_k_index[1486] = 6595;
mem_k_index[1487] = 6598;
mem_k_index[1488] = 6600;
mem_k_index[1489] = 6603;
mem_k_index[1490] = 6605;
mem_k_index[1491] = 6608;
mem_k_index[1492] = 6610;
mem_k_index[1493] = 6613;
mem_k_index[1494] = 6616;
mem_k_index[1495] = 6618;
mem_k_index[1496] = 6621;
mem_k_index[1497] = 6623;
mem_k_index[1498] = 6626;
mem_k_index[1499] = 6628;
mem_k_index[1500] = 6631;
mem_k_index[1501] = 6633;
mem_k_index[1502] = 6636;
mem_k_index[1503] = 6638;
mem_k_index[1504] = 6641;
mem_k_index[1505] = 6643;
mem_k_index[1506] = 6646;
mem_k_index[1507] = 6648;
mem_k_index[1508] = 6651;
mem_k_index[1509] = 6653;
mem_k_index[1510] = 6656;
mem_k_index[1511] = 6658;
mem_k_index[1512] = 6661;
mem_k_index[1513] = 6663;
mem_k_index[1514] = 6666;
mem_k_index[1515] = 6668;
mem_k_index[1516] = 6671;
mem_k_index[1517] = 6673;
mem_k_index[1518] = 6676;
mem_k_index[1519] = 6678;
mem_k_index[1520] = 6681;
mem_k_index[1521] = 6683;
mem_k_index[1522] = 6686;
mem_k_index[1523] = 6688;
mem_k_index[1524] = 6691;
mem_k_index[1525] = 6693;
mem_k_index[1526] = 6696;
mem_k_index[1527] = 6698;
mem_k_index[1528] = 6701;
mem_k_index[1529] = 6703;
mem_k_index[1530] = 6706;
mem_k_index[1531] = 6708;
mem_k_index[1532] = 6711;
mem_k_index[1533] = 6713;
mem_k_index[1534] = 6716;
mem_k_index[1535] = 6718;
mem_k_index[1536] = 7040;
mem_k_index[1537] = 7042;
mem_k_index[1538] = 7045;
mem_k_index[1539] = 7047;
mem_k_index[1540] = 7050;
mem_k_index[1541] = 7052;
mem_k_index[1542] = 7055;
mem_k_index[1543] = 7057;
mem_k_index[1544] = 7060;
mem_k_index[1545] = 7062;
mem_k_index[1546] = 7065;
mem_k_index[1547] = 7067;
mem_k_index[1548] = 7070;
mem_k_index[1549] = 7072;
mem_k_index[1550] = 7075;
mem_k_index[1551] = 7077;
mem_k_index[1552] = 7080;
mem_k_index[1553] = 7082;
mem_k_index[1554] = 7085;
mem_k_index[1555] = 7087;
mem_k_index[1556] = 7090;
mem_k_index[1557] = 7092;
mem_k_index[1558] = 7095;
mem_k_index[1559] = 7097;
mem_k_index[1560] = 7100;
mem_k_index[1561] = 7102;
mem_k_index[1562] = 7105;
mem_k_index[1563] = 7107;
mem_k_index[1564] = 7110;
mem_k_index[1565] = 7112;
mem_k_index[1566] = 7115;
mem_k_index[1567] = 7117;
mem_k_index[1568] = 7120;
mem_k_index[1569] = 7122;
mem_k_index[1570] = 7125;
mem_k_index[1571] = 7127;
mem_k_index[1572] = 7130;
mem_k_index[1573] = 7132;
mem_k_index[1574] = 7135;
mem_k_index[1575] = 7137;
mem_k_index[1576] = 7140;
mem_k_index[1577] = 7142;
mem_k_index[1578] = 7145;
mem_k_index[1579] = 7148;
mem_k_index[1580] = 7150;
mem_k_index[1581] = 7153;
mem_k_index[1582] = 7155;
mem_k_index[1583] = 7158;
mem_k_index[1584] = 7160;
mem_k_index[1585] = 7163;
mem_k_index[1586] = 7165;
mem_k_index[1587] = 7168;
mem_k_index[1588] = 7170;
mem_k_index[1589] = 7173;
mem_k_index[1590] = 7175;
mem_k_index[1591] = 7178;
mem_k_index[1592] = 7180;
mem_k_index[1593] = 7183;
mem_k_index[1594] = 7185;
mem_k_index[1595] = 7188;
mem_k_index[1596] = 7190;
mem_k_index[1597] = 7193;
mem_k_index[1598] = 7195;
mem_k_index[1599] = 7198;
mem_k_index[1600] = 7200;
mem_k_index[1601] = 7203;
mem_k_index[1602] = 7205;
mem_k_index[1603] = 7208;
mem_k_index[1604] = 7210;
mem_k_index[1605] = 7213;
mem_k_index[1606] = 7215;
mem_k_index[1607] = 7218;
mem_k_index[1608] = 7220;
mem_k_index[1609] = 7223;
mem_k_index[1610] = 7225;
mem_k_index[1611] = 7228;
mem_k_index[1612] = 7230;
mem_k_index[1613] = 7233;
mem_k_index[1614] = 7235;
mem_k_index[1615] = 7238;
mem_k_index[1616] = 7240;
mem_k_index[1617] = 7243;
mem_k_index[1618] = 7245;
mem_k_index[1619] = 7248;
mem_k_index[1620] = 7250;
mem_k_index[1621] = 7253;
mem_k_index[1622] = 7256;
mem_k_index[1623] = 7258;
mem_k_index[1624] = 7261;
mem_k_index[1625] = 7263;
mem_k_index[1626] = 7266;
mem_k_index[1627] = 7268;
mem_k_index[1628] = 7271;
mem_k_index[1629] = 7273;
mem_k_index[1630] = 7276;
mem_k_index[1631] = 7278;
mem_k_index[1632] = 7281;
mem_k_index[1633] = 7283;
mem_k_index[1634] = 7286;
mem_k_index[1635] = 7288;
mem_k_index[1636] = 7291;
mem_k_index[1637] = 7293;
mem_k_index[1638] = 7296;
mem_k_index[1639] = 7298;
mem_k_index[1640] = 7301;
mem_k_index[1641] = 7303;
mem_k_index[1642] = 7306;
mem_k_index[1643] = 7308;
mem_k_index[1644] = 7311;
mem_k_index[1645] = 7313;
mem_k_index[1646] = 7316;
mem_k_index[1647] = 7318;
mem_k_index[1648] = 7321;
mem_k_index[1649] = 7323;
mem_k_index[1650] = 7326;
mem_k_index[1651] = 7328;
mem_k_index[1652] = 7331;
mem_k_index[1653] = 7333;
mem_k_index[1654] = 7336;
mem_k_index[1655] = 7338;
mem_k_index[1656] = 7341;
mem_k_index[1657] = 7343;
mem_k_index[1658] = 7346;
mem_k_index[1659] = 7348;
mem_k_index[1660] = 7351;
mem_k_index[1661] = 7353;
mem_k_index[1662] = 7356;
mem_k_index[1663] = 7358;
mem_k_index[1664] = 7680;
mem_k_index[1665] = 7682;
mem_k_index[1666] = 7685;
mem_k_index[1667] = 7687;
mem_k_index[1668] = 7690;
mem_k_index[1669] = 7692;
mem_k_index[1670] = 7695;
mem_k_index[1671] = 7697;
mem_k_index[1672] = 7700;
mem_k_index[1673] = 7702;
mem_k_index[1674] = 7705;
mem_k_index[1675] = 7707;
mem_k_index[1676] = 7710;
mem_k_index[1677] = 7712;
mem_k_index[1678] = 7715;
mem_k_index[1679] = 7717;
mem_k_index[1680] = 7720;
mem_k_index[1681] = 7722;
mem_k_index[1682] = 7725;
mem_k_index[1683] = 7727;
mem_k_index[1684] = 7730;
mem_k_index[1685] = 7732;
mem_k_index[1686] = 7735;
mem_k_index[1687] = 7737;
mem_k_index[1688] = 7740;
mem_k_index[1689] = 7742;
mem_k_index[1690] = 7745;
mem_k_index[1691] = 7747;
mem_k_index[1692] = 7750;
mem_k_index[1693] = 7752;
mem_k_index[1694] = 7755;
mem_k_index[1695] = 7757;
mem_k_index[1696] = 7760;
mem_k_index[1697] = 7762;
mem_k_index[1698] = 7765;
mem_k_index[1699] = 7767;
mem_k_index[1700] = 7770;
mem_k_index[1701] = 7772;
mem_k_index[1702] = 7775;
mem_k_index[1703] = 7777;
mem_k_index[1704] = 7780;
mem_k_index[1705] = 7782;
mem_k_index[1706] = 7785;
mem_k_index[1707] = 7788;
mem_k_index[1708] = 7790;
mem_k_index[1709] = 7793;
mem_k_index[1710] = 7795;
mem_k_index[1711] = 7798;
mem_k_index[1712] = 7800;
mem_k_index[1713] = 7803;
mem_k_index[1714] = 7805;
mem_k_index[1715] = 7808;
mem_k_index[1716] = 7810;
mem_k_index[1717] = 7813;
mem_k_index[1718] = 7815;
mem_k_index[1719] = 7818;
mem_k_index[1720] = 7820;
mem_k_index[1721] = 7823;
mem_k_index[1722] = 7825;
mem_k_index[1723] = 7828;
mem_k_index[1724] = 7830;
mem_k_index[1725] = 7833;
mem_k_index[1726] = 7835;
mem_k_index[1727] = 7838;
mem_k_index[1728] = 7840;
mem_k_index[1729] = 7843;
mem_k_index[1730] = 7845;
mem_k_index[1731] = 7848;
mem_k_index[1732] = 7850;
mem_k_index[1733] = 7853;
mem_k_index[1734] = 7855;
mem_k_index[1735] = 7858;
mem_k_index[1736] = 7860;
mem_k_index[1737] = 7863;
mem_k_index[1738] = 7865;
mem_k_index[1739] = 7868;
mem_k_index[1740] = 7870;
mem_k_index[1741] = 7873;
mem_k_index[1742] = 7875;
mem_k_index[1743] = 7878;
mem_k_index[1744] = 7880;
mem_k_index[1745] = 7883;
mem_k_index[1746] = 7885;
mem_k_index[1747] = 7888;
mem_k_index[1748] = 7890;
mem_k_index[1749] = 7893;
mem_k_index[1750] = 7896;
mem_k_index[1751] = 7898;
mem_k_index[1752] = 7901;
mem_k_index[1753] = 7903;
mem_k_index[1754] = 7906;
mem_k_index[1755] = 7908;
mem_k_index[1756] = 7911;
mem_k_index[1757] = 7913;
mem_k_index[1758] = 7916;
mem_k_index[1759] = 7918;
mem_k_index[1760] = 7921;
mem_k_index[1761] = 7923;
mem_k_index[1762] = 7926;
mem_k_index[1763] = 7928;
mem_k_index[1764] = 7931;
mem_k_index[1765] = 7933;
mem_k_index[1766] = 7936;
mem_k_index[1767] = 7938;
mem_k_index[1768] = 7941;
mem_k_index[1769] = 7943;
mem_k_index[1770] = 7946;
mem_k_index[1771] = 7948;
mem_k_index[1772] = 7951;
mem_k_index[1773] = 7953;
mem_k_index[1774] = 7956;
mem_k_index[1775] = 7958;
mem_k_index[1776] = 7961;
mem_k_index[1777] = 7963;
mem_k_index[1778] = 7966;
mem_k_index[1779] = 7968;
mem_k_index[1780] = 7971;
mem_k_index[1781] = 7973;
mem_k_index[1782] = 7976;
mem_k_index[1783] = 7978;
mem_k_index[1784] = 7981;
mem_k_index[1785] = 7983;
mem_k_index[1786] = 7986;
mem_k_index[1787] = 7988;
mem_k_index[1788] = 7991;
mem_k_index[1789] = 7993;
mem_k_index[1790] = 7996;
mem_k_index[1791] = 7998;
mem_k_index[1792] = 8320;
mem_k_index[1793] = 8322;
mem_k_index[1794] = 8325;
mem_k_index[1795] = 8327;
mem_k_index[1796] = 8330;
mem_k_index[1797] = 8332;
mem_k_index[1798] = 8335;
mem_k_index[1799] = 8337;
mem_k_index[1800] = 8340;
mem_k_index[1801] = 8342;
mem_k_index[1802] = 8345;
mem_k_index[1803] = 8347;
mem_k_index[1804] = 8350;
mem_k_index[1805] = 8352;
mem_k_index[1806] = 8355;
mem_k_index[1807] = 8357;
mem_k_index[1808] = 8360;
mem_k_index[1809] = 8362;
mem_k_index[1810] = 8365;
mem_k_index[1811] = 8367;
mem_k_index[1812] = 8370;
mem_k_index[1813] = 8372;
mem_k_index[1814] = 8375;
mem_k_index[1815] = 8377;
mem_k_index[1816] = 8380;
mem_k_index[1817] = 8382;
mem_k_index[1818] = 8385;
mem_k_index[1819] = 8387;
mem_k_index[1820] = 8390;
mem_k_index[1821] = 8392;
mem_k_index[1822] = 8395;
mem_k_index[1823] = 8397;
mem_k_index[1824] = 8400;
mem_k_index[1825] = 8402;
mem_k_index[1826] = 8405;
mem_k_index[1827] = 8407;
mem_k_index[1828] = 8410;
mem_k_index[1829] = 8412;
mem_k_index[1830] = 8415;
mem_k_index[1831] = 8417;
mem_k_index[1832] = 8420;
mem_k_index[1833] = 8422;
mem_k_index[1834] = 8425;
mem_k_index[1835] = 8428;
mem_k_index[1836] = 8430;
mem_k_index[1837] = 8433;
mem_k_index[1838] = 8435;
mem_k_index[1839] = 8438;
mem_k_index[1840] = 8440;
mem_k_index[1841] = 8443;
mem_k_index[1842] = 8445;
mem_k_index[1843] = 8448;
mem_k_index[1844] = 8450;
mem_k_index[1845] = 8453;
mem_k_index[1846] = 8455;
mem_k_index[1847] = 8458;
mem_k_index[1848] = 8460;
mem_k_index[1849] = 8463;
mem_k_index[1850] = 8465;
mem_k_index[1851] = 8468;
mem_k_index[1852] = 8470;
mem_k_index[1853] = 8473;
mem_k_index[1854] = 8475;
mem_k_index[1855] = 8478;
mem_k_index[1856] = 8480;
mem_k_index[1857] = 8483;
mem_k_index[1858] = 8485;
mem_k_index[1859] = 8488;
mem_k_index[1860] = 8490;
mem_k_index[1861] = 8493;
mem_k_index[1862] = 8495;
mem_k_index[1863] = 8498;
mem_k_index[1864] = 8500;
mem_k_index[1865] = 8503;
mem_k_index[1866] = 8505;
mem_k_index[1867] = 8508;
mem_k_index[1868] = 8510;
mem_k_index[1869] = 8513;
mem_k_index[1870] = 8515;
mem_k_index[1871] = 8518;
mem_k_index[1872] = 8520;
mem_k_index[1873] = 8523;
mem_k_index[1874] = 8525;
mem_k_index[1875] = 8528;
mem_k_index[1876] = 8530;
mem_k_index[1877] = 8533;
mem_k_index[1878] = 8536;
mem_k_index[1879] = 8538;
mem_k_index[1880] = 8541;
mem_k_index[1881] = 8543;
mem_k_index[1882] = 8546;
mem_k_index[1883] = 8548;
mem_k_index[1884] = 8551;
mem_k_index[1885] = 8553;
mem_k_index[1886] = 8556;
mem_k_index[1887] = 8558;
mem_k_index[1888] = 8561;
mem_k_index[1889] = 8563;
mem_k_index[1890] = 8566;
mem_k_index[1891] = 8568;
mem_k_index[1892] = 8571;
mem_k_index[1893] = 8573;
mem_k_index[1894] = 8576;
mem_k_index[1895] = 8578;
mem_k_index[1896] = 8581;
mem_k_index[1897] = 8583;
mem_k_index[1898] = 8586;
mem_k_index[1899] = 8588;
mem_k_index[1900] = 8591;
mem_k_index[1901] = 8593;
mem_k_index[1902] = 8596;
mem_k_index[1903] = 8598;
mem_k_index[1904] = 8601;
mem_k_index[1905] = 8603;
mem_k_index[1906] = 8606;
mem_k_index[1907] = 8608;
mem_k_index[1908] = 8611;
mem_k_index[1909] = 8613;
mem_k_index[1910] = 8616;
mem_k_index[1911] = 8618;
mem_k_index[1912] = 8621;
mem_k_index[1913] = 8623;
mem_k_index[1914] = 8626;
mem_k_index[1915] = 8628;
mem_k_index[1916] = 8631;
mem_k_index[1917] = 8633;
mem_k_index[1918] = 8636;
mem_k_index[1919] = 8638;
mem_k_index[1920] = 8960;
mem_k_index[1921] = 8962;
mem_k_index[1922] = 8965;
mem_k_index[1923] = 8967;
mem_k_index[1924] = 8970;
mem_k_index[1925] = 8972;
mem_k_index[1926] = 8975;
mem_k_index[1927] = 8977;
mem_k_index[1928] = 8980;
mem_k_index[1929] = 8982;
mem_k_index[1930] = 8985;
mem_k_index[1931] = 8987;
mem_k_index[1932] = 8990;
mem_k_index[1933] = 8992;
mem_k_index[1934] = 8995;
mem_k_index[1935] = 8997;
mem_k_index[1936] = 9000;
mem_k_index[1937] = 9002;
mem_k_index[1938] = 9005;
mem_k_index[1939] = 9007;
mem_k_index[1940] = 9010;
mem_k_index[1941] = 9012;
mem_k_index[1942] = 9015;
mem_k_index[1943] = 9017;
mem_k_index[1944] = 9020;
mem_k_index[1945] = 9022;
mem_k_index[1946] = 9025;
mem_k_index[1947] = 9027;
mem_k_index[1948] = 9030;
mem_k_index[1949] = 9032;
mem_k_index[1950] = 9035;
mem_k_index[1951] = 9037;
mem_k_index[1952] = 9040;
mem_k_index[1953] = 9042;
mem_k_index[1954] = 9045;
mem_k_index[1955] = 9047;
mem_k_index[1956] = 9050;
mem_k_index[1957] = 9052;
mem_k_index[1958] = 9055;
mem_k_index[1959] = 9057;
mem_k_index[1960] = 9060;
mem_k_index[1961] = 9062;
mem_k_index[1962] = 9065;
mem_k_index[1963] = 9068;
mem_k_index[1964] = 9070;
mem_k_index[1965] = 9073;
mem_k_index[1966] = 9075;
mem_k_index[1967] = 9078;
mem_k_index[1968] = 9080;
mem_k_index[1969] = 9083;
mem_k_index[1970] = 9085;
mem_k_index[1971] = 9088;
mem_k_index[1972] = 9090;
mem_k_index[1973] = 9093;
mem_k_index[1974] = 9095;
mem_k_index[1975] = 9098;
mem_k_index[1976] = 9100;
mem_k_index[1977] = 9103;
mem_k_index[1978] = 9105;
mem_k_index[1979] = 9108;
mem_k_index[1980] = 9110;
mem_k_index[1981] = 9113;
mem_k_index[1982] = 9115;
mem_k_index[1983] = 9118;
mem_k_index[1984] = 9120;
mem_k_index[1985] = 9123;
mem_k_index[1986] = 9125;
mem_k_index[1987] = 9128;
mem_k_index[1988] = 9130;
mem_k_index[1989] = 9133;
mem_k_index[1990] = 9135;
mem_k_index[1991] = 9138;
mem_k_index[1992] = 9140;
mem_k_index[1993] = 9143;
mem_k_index[1994] = 9145;
mem_k_index[1995] = 9148;
mem_k_index[1996] = 9150;
mem_k_index[1997] = 9153;
mem_k_index[1998] = 9155;
mem_k_index[1999] = 9158;
mem_k_index[2000] = 9160;
mem_k_index[2001] = 9163;
mem_k_index[2002] = 9165;
mem_k_index[2003] = 9168;
mem_k_index[2004] = 9170;
mem_k_index[2005] = 9173;
mem_k_index[2006] = 9176;
mem_k_index[2007] = 9178;
mem_k_index[2008] = 9181;
mem_k_index[2009] = 9183;
mem_k_index[2010] = 9186;
mem_k_index[2011] = 9188;
mem_k_index[2012] = 9191;
mem_k_index[2013] = 9193;
mem_k_index[2014] = 9196;
mem_k_index[2015] = 9198;
mem_k_index[2016] = 9201;
mem_k_index[2017] = 9203;
mem_k_index[2018] = 9206;
mem_k_index[2019] = 9208;
mem_k_index[2020] = 9211;
mem_k_index[2021] = 9213;
mem_k_index[2022] = 9216;
mem_k_index[2023] = 9218;
mem_k_index[2024] = 9221;
mem_k_index[2025] = 9223;
mem_k_index[2026] = 9226;
mem_k_index[2027] = 9228;
mem_k_index[2028] = 9231;
mem_k_index[2029] = 9233;
mem_k_index[2030] = 9236;
mem_k_index[2031] = 9238;
mem_k_index[2032] = 9241;
mem_k_index[2033] = 9243;
mem_k_index[2034] = 9246;
mem_k_index[2035] = 9248;
mem_k_index[2036] = 9251;
mem_k_index[2037] = 9253;
mem_k_index[2038] = 9256;
mem_k_index[2039] = 9258;
mem_k_index[2040] = 9261;
mem_k_index[2041] = 9263;
mem_k_index[2042] = 9266;
mem_k_index[2043] = 9268;
mem_k_index[2044] = 9271;
mem_k_index[2045] = 9273;
mem_k_index[2046] = 9276;
mem_k_index[2047] = 9278;
mem_k_index[2048] = 9600;
mem_k_index[2049] = 9602;
mem_k_index[2050] = 9605;
mem_k_index[2051] = 9607;
mem_k_index[2052] = 9610;
mem_k_index[2053] = 9612;
mem_k_index[2054] = 9615;
mem_k_index[2055] = 9617;
mem_k_index[2056] = 9620;
mem_k_index[2057] = 9622;
mem_k_index[2058] = 9625;
mem_k_index[2059] = 9627;
mem_k_index[2060] = 9630;
mem_k_index[2061] = 9632;
mem_k_index[2062] = 9635;
mem_k_index[2063] = 9637;
mem_k_index[2064] = 9640;
mem_k_index[2065] = 9642;
mem_k_index[2066] = 9645;
mem_k_index[2067] = 9647;
mem_k_index[2068] = 9650;
mem_k_index[2069] = 9652;
mem_k_index[2070] = 9655;
mem_k_index[2071] = 9657;
mem_k_index[2072] = 9660;
mem_k_index[2073] = 9662;
mem_k_index[2074] = 9665;
mem_k_index[2075] = 9667;
mem_k_index[2076] = 9670;
mem_k_index[2077] = 9672;
mem_k_index[2078] = 9675;
mem_k_index[2079] = 9677;
mem_k_index[2080] = 9680;
mem_k_index[2081] = 9682;
mem_k_index[2082] = 9685;
mem_k_index[2083] = 9687;
mem_k_index[2084] = 9690;
mem_k_index[2085] = 9692;
mem_k_index[2086] = 9695;
mem_k_index[2087] = 9697;
mem_k_index[2088] = 9700;
mem_k_index[2089] = 9702;
mem_k_index[2090] = 9705;
mem_k_index[2091] = 9708;
mem_k_index[2092] = 9710;
mem_k_index[2093] = 9713;
mem_k_index[2094] = 9715;
mem_k_index[2095] = 9718;
mem_k_index[2096] = 9720;
mem_k_index[2097] = 9723;
mem_k_index[2098] = 9725;
mem_k_index[2099] = 9728;
mem_k_index[2100] = 9730;
mem_k_index[2101] = 9733;
mem_k_index[2102] = 9735;
mem_k_index[2103] = 9738;
mem_k_index[2104] = 9740;
mem_k_index[2105] = 9743;
mem_k_index[2106] = 9745;
mem_k_index[2107] = 9748;
mem_k_index[2108] = 9750;
mem_k_index[2109] = 9753;
mem_k_index[2110] = 9755;
mem_k_index[2111] = 9758;
mem_k_index[2112] = 9760;
mem_k_index[2113] = 9763;
mem_k_index[2114] = 9765;
mem_k_index[2115] = 9768;
mem_k_index[2116] = 9770;
mem_k_index[2117] = 9773;
mem_k_index[2118] = 9775;
mem_k_index[2119] = 9778;
mem_k_index[2120] = 9780;
mem_k_index[2121] = 9783;
mem_k_index[2122] = 9785;
mem_k_index[2123] = 9788;
mem_k_index[2124] = 9790;
mem_k_index[2125] = 9793;
mem_k_index[2126] = 9795;
mem_k_index[2127] = 9798;
mem_k_index[2128] = 9800;
mem_k_index[2129] = 9803;
mem_k_index[2130] = 9805;
mem_k_index[2131] = 9808;
mem_k_index[2132] = 9810;
mem_k_index[2133] = 9813;
mem_k_index[2134] = 9816;
mem_k_index[2135] = 9818;
mem_k_index[2136] = 9821;
mem_k_index[2137] = 9823;
mem_k_index[2138] = 9826;
mem_k_index[2139] = 9828;
mem_k_index[2140] = 9831;
mem_k_index[2141] = 9833;
mem_k_index[2142] = 9836;
mem_k_index[2143] = 9838;
mem_k_index[2144] = 9841;
mem_k_index[2145] = 9843;
mem_k_index[2146] = 9846;
mem_k_index[2147] = 9848;
mem_k_index[2148] = 9851;
mem_k_index[2149] = 9853;
mem_k_index[2150] = 9856;
mem_k_index[2151] = 9858;
mem_k_index[2152] = 9861;
mem_k_index[2153] = 9863;
mem_k_index[2154] = 9866;
mem_k_index[2155] = 9868;
mem_k_index[2156] = 9871;
mem_k_index[2157] = 9873;
mem_k_index[2158] = 9876;
mem_k_index[2159] = 9878;
mem_k_index[2160] = 9881;
mem_k_index[2161] = 9883;
mem_k_index[2162] = 9886;
mem_k_index[2163] = 9888;
mem_k_index[2164] = 9891;
mem_k_index[2165] = 9893;
mem_k_index[2166] = 9896;
mem_k_index[2167] = 9898;
mem_k_index[2168] = 9901;
mem_k_index[2169] = 9903;
mem_k_index[2170] = 9906;
mem_k_index[2171] = 9908;
mem_k_index[2172] = 9911;
mem_k_index[2173] = 9913;
mem_k_index[2174] = 9916;
mem_k_index[2175] = 9918;
mem_k_index[2176] = 9920;
mem_k_index[2177] = 9922;
mem_k_index[2178] = 9925;
mem_k_index[2179] = 9927;
mem_k_index[2180] = 9930;
mem_k_index[2181] = 9932;
mem_k_index[2182] = 9935;
mem_k_index[2183] = 9937;
mem_k_index[2184] = 9940;
mem_k_index[2185] = 9942;
mem_k_index[2186] = 9945;
mem_k_index[2187] = 9947;
mem_k_index[2188] = 9950;
mem_k_index[2189] = 9952;
mem_k_index[2190] = 9955;
mem_k_index[2191] = 9957;
mem_k_index[2192] = 9960;
mem_k_index[2193] = 9962;
mem_k_index[2194] = 9965;
mem_k_index[2195] = 9967;
mem_k_index[2196] = 9970;
mem_k_index[2197] = 9972;
mem_k_index[2198] = 9975;
mem_k_index[2199] = 9977;
mem_k_index[2200] = 9980;
mem_k_index[2201] = 9982;
mem_k_index[2202] = 9985;
mem_k_index[2203] = 9987;
mem_k_index[2204] = 9990;
mem_k_index[2205] = 9992;
mem_k_index[2206] = 9995;
mem_k_index[2207] = 9997;
mem_k_index[2208] = 10000;
mem_k_index[2209] = 10002;
mem_k_index[2210] = 10005;
mem_k_index[2211] = 10007;
mem_k_index[2212] = 10010;
mem_k_index[2213] = 10012;
mem_k_index[2214] = 10015;
mem_k_index[2215] = 10017;
mem_k_index[2216] = 10020;
mem_k_index[2217] = 10022;
mem_k_index[2218] = 10025;
mem_k_index[2219] = 10028;
mem_k_index[2220] = 10030;
mem_k_index[2221] = 10033;
mem_k_index[2222] = 10035;
mem_k_index[2223] = 10038;
mem_k_index[2224] = 10040;
mem_k_index[2225] = 10043;
mem_k_index[2226] = 10045;
mem_k_index[2227] = 10048;
mem_k_index[2228] = 10050;
mem_k_index[2229] = 10053;
mem_k_index[2230] = 10055;
mem_k_index[2231] = 10058;
mem_k_index[2232] = 10060;
mem_k_index[2233] = 10063;
mem_k_index[2234] = 10065;
mem_k_index[2235] = 10068;
mem_k_index[2236] = 10070;
mem_k_index[2237] = 10073;
mem_k_index[2238] = 10075;
mem_k_index[2239] = 10078;
mem_k_index[2240] = 10080;
mem_k_index[2241] = 10083;
mem_k_index[2242] = 10085;
mem_k_index[2243] = 10088;
mem_k_index[2244] = 10090;
mem_k_index[2245] = 10093;
mem_k_index[2246] = 10095;
mem_k_index[2247] = 10098;
mem_k_index[2248] = 10100;
mem_k_index[2249] = 10103;
mem_k_index[2250] = 10105;
mem_k_index[2251] = 10108;
mem_k_index[2252] = 10110;
mem_k_index[2253] = 10113;
mem_k_index[2254] = 10115;
mem_k_index[2255] = 10118;
mem_k_index[2256] = 10120;
mem_k_index[2257] = 10123;
mem_k_index[2258] = 10125;
mem_k_index[2259] = 10128;
mem_k_index[2260] = 10130;
mem_k_index[2261] = 10133;
mem_k_index[2262] = 10136;
mem_k_index[2263] = 10138;
mem_k_index[2264] = 10141;
mem_k_index[2265] = 10143;
mem_k_index[2266] = 10146;
mem_k_index[2267] = 10148;
mem_k_index[2268] = 10151;
mem_k_index[2269] = 10153;
mem_k_index[2270] = 10156;
mem_k_index[2271] = 10158;
mem_k_index[2272] = 10161;
mem_k_index[2273] = 10163;
mem_k_index[2274] = 10166;
mem_k_index[2275] = 10168;
mem_k_index[2276] = 10171;
mem_k_index[2277] = 10173;
mem_k_index[2278] = 10176;
mem_k_index[2279] = 10178;
mem_k_index[2280] = 10181;
mem_k_index[2281] = 10183;
mem_k_index[2282] = 10186;
mem_k_index[2283] = 10188;
mem_k_index[2284] = 10191;
mem_k_index[2285] = 10193;
mem_k_index[2286] = 10196;
mem_k_index[2287] = 10198;
mem_k_index[2288] = 10201;
mem_k_index[2289] = 10203;
mem_k_index[2290] = 10206;
mem_k_index[2291] = 10208;
mem_k_index[2292] = 10211;
mem_k_index[2293] = 10213;
mem_k_index[2294] = 10216;
mem_k_index[2295] = 10218;
mem_k_index[2296] = 10221;
mem_k_index[2297] = 10223;
mem_k_index[2298] = 10226;
mem_k_index[2299] = 10228;
mem_k_index[2300] = 10231;
mem_k_index[2301] = 10233;
mem_k_index[2302] = 10236;
mem_k_index[2303] = 10238;
mem_k_index[2304] = 10560;
mem_k_index[2305] = 10562;
mem_k_index[2306] = 10565;
mem_k_index[2307] = 10567;
mem_k_index[2308] = 10570;
mem_k_index[2309] = 10572;
mem_k_index[2310] = 10575;
mem_k_index[2311] = 10577;
mem_k_index[2312] = 10580;
mem_k_index[2313] = 10582;
mem_k_index[2314] = 10585;
mem_k_index[2315] = 10587;
mem_k_index[2316] = 10590;
mem_k_index[2317] = 10592;
mem_k_index[2318] = 10595;
mem_k_index[2319] = 10597;
mem_k_index[2320] = 10600;
mem_k_index[2321] = 10602;
mem_k_index[2322] = 10605;
mem_k_index[2323] = 10607;
mem_k_index[2324] = 10610;
mem_k_index[2325] = 10612;
mem_k_index[2326] = 10615;
mem_k_index[2327] = 10617;
mem_k_index[2328] = 10620;
mem_k_index[2329] = 10622;
mem_k_index[2330] = 10625;
mem_k_index[2331] = 10627;
mem_k_index[2332] = 10630;
mem_k_index[2333] = 10632;
mem_k_index[2334] = 10635;
mem_k_index[2335] = 10637;
mem_k_index[2336] = 10640;
mem_k_index[2337] = 10642;
mem_k_index[2338] = 10645;
mem_k_index[2339] = 10647;
mem_k_index[2340] = 10650;
mem_k_index[2341] = 10652;
mem_k_index[2342] = 10655;
mem_k_index[2343] = 10657;
mem_k_index[2344] = 10660;
mem_k_index[2345] = 10662;
mem_k_index[2346] = 10665;
mem_k_index[2347] = 10668;
mem_k_index[2348] = 10670;
mem_k_index[2349] = 10673;
mem_k_index[2350] = 10675;
mem_k_index[2351] = 10678;
mem_k_index[2352] = 10680;
mem_k_index[2353] = 10683;
mem_k_index[2354] = 10685;
mem_k_index[2355] = 10688;
mem_k_index[2356] = 10690;
mem_k_index[2357] = 10693;
mem_k_index[2358] = 10695;
mem_k_index[2359] = 10698;
mem_k_index[2360] = 10700;
mem_k_index[2361] = 10703;
mem_k_index[2362] = 10705;
mem_k_index[2363] = 10708;
mem_k_index[2364] = 10710;
mem_k_index[2365] = 10713;
mem_k_index[2366] = 10715;
mem_k_index[2367] = 10718;
mem_k_index[2368] = 10720;
mem_k_index[2369] = 10723;
mem_k_index[2370] = 10725;
mem_k_index[2371] = 10728;
mem_k_index[2372] = 10730;
mem_k_index[2373] = 10733;
mem_k_index[2374] = 10735;
mem_k_index[2375] = 10738;
mem_k_index[2376] = 10740;
mem_k_index[2377] = 10743;
mem_k_index[2378] = 10745;
mem_k_index[2379] = 10748;
mem_k_index[2380] = 10750;
mem_k_index[2381] = 10753;
mem_k_index[2382] = 10755;
mem_k_index[2383] = 10758;
mem_k_index[2384] = 10760;
mem_k_index[2385] = 10763;
mem_k_index[2386] = 10765;
mem_k_index[2387] = 10768;
mem_k_index[2388] = 10770;
mem_k_index[2389] = 10773;
mem_k_index[2390] = 10776;
mem_k_index[2391] = 10778;
mem_k_index[2392] = 10781;
mem_k_index[2393] = 10783;
mem_k_index[2394] = 10786;
mem_k_index[2395] = 10788;
mem_k_index[2396] = 10791;
mem_k_index[2397] = 10793;
mem_k_index[2398] = 10796;
mem_k_index[2399] = 10798;
mem_k_index[2400] = 10801;
mem_k_index[2401] = 10803;
mem_k_index[2402] = 10806;
mem_k_index[2403] = 10808;
mem_k_index[2404] = 10811;
mem_k_index[2405] = 10813;
mem_k_index[2406] = 10816;
mem_k_index[2407] = 10818;
mem_k_index[2408] = 10821;
mem_k_index[2409] = 10823;
mem_k_index[2410] = 10826;
mem_k_index[2411] = 10828;
mem_k_index[2412] = 10831;
mem_k_index[2413] = 10833;
mem_k_index[2414] = 10836;
mem_k_index[2415] = 10838;
mem_k_index[2416] = 10841;
mem_k_index[2417] = 10843;
mem_k_index[2418] = 10846;
mem_k_index[2419] = 10848;
mem_k_index[2420] = 10851;
mem_k_index[2421] = 10853;
mem_k_index[2422] = 10856;
mem_k_index[2423] = 10858;
mem_k_index[2424] = 10861;
mem_k_index[2425] = 10863;
mem_k_index[2426] = 10866;
mem_k_index[2427] = 10868;
mem_k_index[2428] = 10871;
mem_k_index[2429] = 10873;
mem_k_index[2430] = 10876;
mem_k_index[2431] = 10878;
mem_k_index[2432] = 11200;
mem_k_index[2433] = 11202;
mem_k_index[2434] = 11205;
mem_k_index[2435] = 11207;
mem_k_index[2436] = 11210;
mem_k_index[2437] = 11212;
mem_k_index[2438] = 11215;
mem_k_index[2439] = 11217;
mem_k_index[2440] = 11220;
mem_k_index[2441] = 11222;
mem_k_index[2442] = 11225;
mem_k_index[2443] = 11227;
mem_k_index[2444] = 11230;
mem_k_index[2445] = 11232;
mem_k_index[2446] = 11235;
mem_k_index[2447] = 11237;
mem_k_index[2448] = 11240;
mem_k_index[2449] = 11242;
mem_k_index[2450] = 11245;
mem_k_index[2451] = 11247;
mem_k_index[2452] = 11250;
mem_k_index[2453] = 11252;
mem_k_index[2454] = 11255;
mem_k_index[2455] = 11257;
mem_k_index[2456] = 11260;
mem_k_index[2457] = 11262;
mem_k_index[2458] = 11265;
mem_k_index[2459] = 11267;
mem_k_index[2460] = 11270;
mem_k_index[2461] = 11272;
mem_k_index[2462] = 11275;
mem_k_index[2463] = 11277;
mem_k_index[2464] = 11280;
mem_k_index[2465] = 11282;
mem_k_index[2466] = 11285;
mem_k_index[2467] = 11287;
mem_k_index[2468] = 11290;
mem_k_index[2469] = 11292;
mem_k_index[2470] = 11295;
mem_k_index[2471] = 11297;
mem_k_index[2472] = 11300;
mem_k_index[2473] = 11302;
mem_k_index[2474] = 11305;
mem_k_index[2475] = 11308;
mem_k_index[2476] = 11310;
mem_k_index[2477] = 11313;
mem_k_index[2478] = 11315;
mem_k_index[2479] = 11318;
mem_k_index[2480] = 11320;
mem_k_index[2481] = 11323;
mem_k_index[2482] = 11325;
mem_k_index[2483] = 11328;
mem_k_index[2484] = 11330;
mem_k_index[2485] = 11333;
mem_k_index[2486] = 11335;
mem_k_index[2487] = 11338;
mem_k_index[2488] = 11340;
mem_k_index[2489] = 11343;
mem_k_index[2490] = 11345;
mem_k_index[2491] = 11348;
mem_k_index[2492] = 11350;
mem_k_index[2493] = 11353;
mem_k_index[2494] = 11355;
mem_k_index[2495] = 11358;
mem_k_index[2496] = 11360;
mem_k_index[2497] = 11363;
mem_k_index[2498] = 11365;
mem_k_index[2499] = 11368;
mem_k_index[2500] = 11370;
mem_k_index[2501] = 11373;
mem_k_index[2502] = 11375;
mem_k_index[2503] = 11378;
mem_k_index[2504] = 11380;
mem_k_index[2505] = 11383;
mem_k_index[2506] = 11385;
mem_k_index[2507] = 11388;
mem_k_index[2508] = 11390;
mem_k_index[2509] = 11393;
mem_k_index[2510] = 11395;
mem_k_index[2511] = 11398;
mem_k_index[2512] = 11400;
mem_k_index[2513] = 11403;
mem_k_index[2514] = 11405;
mem_k_index[2515] = 11408;
mem_k_index[2516] = 11410;
mem_k_index[2517] = 11413;
mem_k_index[2518] = 11416;
mem_k_index[2519] = 11418;
mem_k_index[2520] = 11421;
mem_k_index[2521] = 11423;
mem_k_index[2522] = 11426;
mem_k_index[2523] = 11428;
mem_k_index[2524] = 11431;
mem_k_index[2525] = 11433;
mem_k_index[2526] = 11436;
mem_k_index[2527] = 11438;
mem_k_index[2528] = 11441;
mem_k_index[2529] = 11443;
mem_k_index[2530] = 11446;
mem_k_index[2531] = 11448;
mem_k_index[2532] = 11451;
mem_k_index[2533] = 11453;
mem_k_index[2534] = 11456;
mem_k_index[2535] = 11458;
mem_k_index[2536] = 11461;
mem_k_index[2537] = 11463;
mem_k_index[2538] = 11466;
mem_k_index[2539] = 11468;
mem_k_index[2540] = 11471;
mem_k_index[2541] = 11473;
mem_k_index[2542] = 11476;
mem_k_index[2543] = 11478;
mem_k_index[2544] = 11481;
mem_k_index[2545] = 11483;
mem_k_index[2546] = 11486;
mem_k_index[2547] = 11488;
mem_k_index[2548] = 11491;
mem_k_index[2549] = 11493;
mem_k_index[2550] = 11496;
mem_k_index[2551] = 11498;
mem_k_index[2552] = 11501;
mem_k_index[2553] = 11503;
mem_k_index[2554] = 11506;
mem_k_index[2555] = 11508;
mem_k_index[2556] = 11511;
mem_k_index[2557] = 11513;
mem_k_index[2558] = 11516;
mem_k_index[2559] = 11518;
mem_k_index[2560] = 11840;
mem_k_index[2561] = 11842;
mem_k_index[2562] = 11845;
mem_k_index[2563] = 11847;
mem_k_index[2564] = 11850;
mem_k_index[2565] = 11852;
mem_k_index[2566] = 11855;
mem_k_index[2567] = 11857;
mem_k_index[2568] = 11860;
mem_k_index[2569] = 11862;
mem_k_index[2570] = 11865;
mem_k_index[2571] = 11867;
mem_k_index[2572] = 11870;
mem_k_index[2573] = 11872;
mem_k_index[2574] = 11875;
mem_k_index[2575] = 11877;
mem_k_index[2576] = 11880;
mem_k_index[2577] = 11882;
mem_k_index[2578] = 11885;
mem_k_index[2579] = 11887;
mem_k_index[2580] = 11890;
mem_k_index[2581] = 11892;
mem_k_index[2582] = 11895;
mem_k_index[2583] = 11897;
mem_k_index[2584] = 11900;
mem_k_index[2585] = 11902;
mem_k_index[2586] = 11905;
mem_k_index[2587] = 11907;
mem_k_index[2588] = 11910;
mem_k_index[2589] = 11912;
mem_k_index[2590] = 11915;
mem_k_index[2591] = 11917;
mem_k_index[2592] = 11920;
mem_k_index[2593] = 11922;
mem_k_index[2594] = 11925;
mem_k_index[2595] = 11927;
mem_k_index[2596] = 11930;
mem_k_index[2597] = 11932;
mem_k_index[2598] = 11935;
mem_k_index[2599] = 11937;
mem_k_index[2600] = 11940;
mem_k_index[2601] = 11942;
mem_k_index[2602] = 11945;
mem_k_index[2603] = 11948;
mem_k_index[2604] = 11950;
mem_k_index[2605] = 11953;
mem_k_index[2606] = 11955;
mem_k_index[2607] = 11958;
mem_k_index[2608] = 11960;
mem_k_index[2609] = 11963;
mem_k_index[2610] = 11965;
mem_k_index[2611] = 11968;
mem_k_index[2612] = 11970;
mem_k_index[2613] = 11973;
mem_k_index[2614] = 11975;
mem_k_index[2615] = 11978;
mem_k_index[2616] = 11980;
mem_k_index[2617] = 11983;
mem_k_index[2618] = 11985;
mem_k_index[2619] = 11988;
mem_k_index[2620] = 11990;
mem_k_index[2621] = 11993;
mem_k_index[2622] = 11995;
mem_k_index[2623] = 11998;
mem_k_index[2624] = 12000;
mem_k_index[2625] = 12003;
mem_k_index[2626] = 12005;
mem_k_index[2627] = 12008;
mem_k_index[2628] = 12010;
mem_k_index[2629] = 12013;
mem_k_index[2630] = 12015;
mem_k_index[2631] = 12018;
mem_k_index[2632] = 12020;
mem_k_index[2633] = 12023;
mem_k_index[2634] = 12025;
mem_k_index[2635] = 12028;
mem_k_index[2636] = 12030;
mem_k_index[2637] = 12033;
mem_k_index[2638] = 12035;
mem_k_index[2639] = 12038;
mem_k_index[2640] = 12040;
mem_k_index[2641] = 12043;
mem_k_index[2642] = 12045;
mem_k_index[2643] = 12048;
mem_k_index[2644] = 12050;
mem_k_index[2645] = 12053;
mem_k_index[2646] = 12056;
mem_k_index[2647] = 12058;
mem_k_index[2648] = 12061;
mem_k_index[2649] = 12063;
mem_k_index[2650] = 12066;
mem_k_index[2651] = 12068;
mem_k_index[2652] = 12071;
mem_k_index[2653] = 12073;
mem_k_index[2654] = 12076;
mem_k_index[2655] = 12078;
mem_k_index[2656] = 12081;
mem_k_index[2657] = 12083;
mem_k_index[2658] = 12086;
mem_k_index[2659] = 12088;
mem_k_index[2660] = 12091;
mem_k_index[2661] = 12093;
mem_k_index[2662] = 12096;
mem_k_index[2663] = 12098;
mem_k_index[2664] = 12101;
mem_k_index[2665] = 12103;
mem_k_index[2666] = 12106;
mem_k_index[2667] = 12108;
mem_k_index[2668] = 12111;
mem_k_index[2669] = 12113;
mem_k_index[2670] = 12116;
mem_k_index[2671] = 12118;
mem_k_index[2672] = 12121;
mem_k_index[2673] = 12123;
mem_k_index[2674] = 12126;
mem_k_index[2675] = 12128;
mem_k_index[2676] = 12131;
mem_k_index[2677] = 12133;
mem_k_index[2678] = 12136;
mem_k_index[2679] = 12138;
mem_k_index[2680] = 12141;
mem_k_index[2681] = 12143;
mem_k_index[2682] = 12146;
mem_k_index[2683] = 12148;
mem_k_index[2684] = 12151;
mem_k_index[2685] = 12153;
mem_k_index[2686] = 12156;
mem_k_index[2687] = 12158;
mem_k_index[2688] = 12480;
mem_k_index[2689] = 12482;
mem_k_index[2690] = 12485;
mem_k_index[2691] = 12487;
mem_k_index[2692] = 12490;
mem_k_index[2693] = 12492;
mem_k_index[2694] = 12495;
mem_k_index[2695] = 12497;
mem_k_index[2696] = 12500;
mem_k_index[2697] = 12502;
mem_k_index[2698] = 12505;
mem_k_index[2699] = 12507;
mem_k_index[2700] = 12510;
mem_k_index[2701] = 12512;
mem_k_index[2702] = 12515;
mem_k_index[2703] = 12517;
mem_k_index[2704] = 12520;
mem_k_index[2705] = 12522;
mem_k_index[2706] = 12525;
mem_k_index[2707] = 12527;
mem_k_index[2708] = 12530;
mem_k_index[2709] = 12532;
mem_k_index[2710] = 12535;
mem_k_index[2711] = 12537;
mem_k_index[2712] = 12540;
mem_k_index[2713] = 12542;
mem_k_index[2714] = 12545;
mem_k_index[2715] = 12547;
mem_k_index[2716] = 12550;
mem_k_index[2717] = 12552;
mem_k_index[2718] = 12555;
mem_k_index[2719] = 12557;
mem_k_index[2720] = 12560;
mem_k_index[2721] = 12562;
mem_k_index[2722] = 12565;
mem_k_index[2723] = 12567;
mem_k_index[2724] = 12570;
mem_k_index[2725] = 12572;
mem_k_index[2726] = 12575;
mem_k_index[2727] = 12577;
mem_k_index[2728] = 12580;
mem_k_index[2729] = 12582;
mem_k_index[2730] = 12585;
mem_k_index[2731] = 12588;
mem_k_index[2732] = 12590;
mem_k_index[2733] = 12593;
mem_k_index[2734] = 12595;
mem_k_index[2735] = 12598;
mem_k_index[2736] = 12600;
mem_k_index[2737] = 12603;
mem_k_index[2738] = 12605;
mem_k_index[2739] = 12608;
mem_k_index[2740] = 12610;
mem_k_index[2741] = 12613;
mem_k_index[2742] = 12615;
mem_k_index[2743] = 12618;
mem_k_index[2744] = 12620;
mem_k_index[2745] = 12623;
mem_k_index[2746] = 12625;
mem_k_index[2747] = 12628;
mem_k_index[2748] = 12630;
mem_k_index[2749] = 12633;
mem_k_index[2750] = 12635;
mem_k_index[2751] = 12638;
mem_k_index[2752] = 12640;
mem_k_index[2753] = 12643;
mem_k_index[2754] = 12645;
mem_k_index[2755] = 12648;
mem_k_index[2756] = 12650;
mem_k_index[2757] = 12653;
mem_k_index[2758] = 12655;
mem_k_index[2759] = 12658;
mem_k_index[2760] = 12660;
mem_k_index[2761] = 12663;
mem_k_index[2762] = 12665;
mem_k_index[2763] = 12668;
mem_k_index[2764] = 12670;
mem_k_index[2765] = 12673;
mem_k_index[2766] = 12675;
mem_k_index[2767] = 12678;
mem_k_index[2768] = 12680;
mem_k_index[2769] = 12683;
mem_k_index[2770] = 12685;
mem_k_index[2771] = 12688;
mem_k_index[2772] = 12690;
mem_k_index[2773] = 12693;
mem_k_index[2774] = 12696;
mem_k_index[2775] = 12698;
mem_k_index[2776] = 12701;
mem_k_index[2777] = 12703;
mem_k_index[2778] = 12706;
mem_k_index[2779] = 12708;
mem_k_index[2780] = 12711;
mem_k_index[2781] = 12713;
mem_k_index[2782] = 12716;
mem_k_index[2783] = 12718;
mem_k_index[2784] = 12721;
mem_k_index[2785] = 12723;
mem_k_index[2786] = 12726;
mem_k_index[2787] = 12728;
mem_k_index[2788] = 12731;
mem_k_index[2789] = 12733;
mem_k_index[2790] = 12736;
mem_k_index[2791] = 12738;
mem_k_index[2792] = 12741;
mem_k_index[2793] = 12743;
mem_k_index[2794] = 12746;
mem_k_index[2795] = 12748;
mem_k_index[2796] = 12751;
mem_k_index[2797] = 12753;
mem_k_index[2798] = 12756;
mem_k_index[2799] = 12758;
mem_k_index[2800] = 12761;
mem_k_index[2801] = 12763;
mem_k_index[2802] = 12766;
mem_k_index[2803] = 12768;
mem_k_index[2804] = 12771;
mem_k_index[2805] = 12773;
mem_k_index[2806] = 12776;
mem_k_index[2807] = 12778;
mem_k_index[2808] = 12781;
mem_k_index[2809] = 12783;
mem_k_index[2810] = 12786;
mem_k_index[2811] = 12788;
mem_k_index[2812] = 12791;
mem_k_index[2813] = 12793;
mem_k_index[2814] = 12796;
mem_k_index[2815] = 12798;
mem_k_index[2816] = 13120;
mem_k_index[2817] = 13122;
mem_k_index[2818] = 13125;
mem_k_index[2819] = 13127;
mem_k_index[2820] = 13130;
mem_k_index[2821] = 13132;
mem_k_index[2822] = 13135;
mem_k_index[2823] = 13137;
mem_k_index[2824] = 13140;
mem_k_index[2825] = 13142;
mem_k_index[2826] = 13145;
mem_k_index[2827] = 13147;
mem_k_index[2828] = 13150;
mem_k_index[2829] = 13152;
mem_k_index[2830] = 13155;
mem_k_index[2831] = 13157;
mem_k_index[2832] = 13160;
mem_k_index[2833] = 13162;
mem_k_index[2834] = 13165;
mem_k_index[2835] = 13167;
mem_k_index[2836] = 13170;
mem_k_index[2837] = 13172;
mem_k_index[2838] = 13175;
mem_k_index[2839] = 13177;
mem_k_index[2840] = 13180;
mem_k_index[2841] = 13182;
mem_k_index[2842] = 13185;
mem_k_index[2843] = 13187;
mem_k_index[2844] = 13190;
mem_k_index[2845] = 13192;
mem_k_index[2846] = 13195;
mem_k_index[2847] = 13197;
mem_k_index[2848] = 13200;
mem_k_index[2849] = 13202;
mem_k_index[2850] = 13205;
mem_k_index[2851] = 13207;
mem_k_index[2852] = 13210;
mem_k_index[2853] = 13212;
mem_k_index[2854] = 13215;
mem_k_index[2855] = 13217;
mem_k_index[2856] = 13220;
mem_k_index[2857] = 13222;
mem_k_index[2858] = 13225;
mem_k_index[2859] = 13228;
mem_k_index[2860] = 13230;
mem_k_index[2861] = 13233;
mem_k_index[2862] = 13235;
mem_k_index[2863] = 13238;
mem_k_index[2864] = 13240;
mem_k_index[2865] = 13243;
mem_k_index[2866] = 13245;
mem_k_index[2867] = 13248;
mem_k_index[2868] = 13250;
mem_k_index[2869] = 13253;
mem_k_index[2870] = 13255;
mem_k_index[2871] = 13258;
mem_k_index[2872] = 13260;
mem_k_index[2873] = 13263;
mem_k_index[2874] = 13265;
mem_k_index[2875] = 13268;
mem_k_index[2876] = 13270;
mem_k_index[2877] = 13273;
mem_k_index[2878] = 13275;
mem_k_index[2879] = 13278;
mem_k_index[2880] = 13280;
mem_k_index[2881] = 13283;
mem_k_index[2882] = 13285;
mem_k_index[2883] = 13288;
mem_k_index[2884] = 13290;
mem_k_index[2885] = 13293;
mem_k_index[2886] = 13295;
mem_k_index[2887] = 13298;
mem_k_index[2888] = 13300;
mem_k_index[2889] = 13303;
mem_k_index[2890] = 13305;
mem_k_index[2891] = 13308;
mem_k_index[2892] = 13310;
mem_k_index[2893] = 13313;
mem_k_index[2894] = 13315;
mem_k_index[2895] = 13318;
mem_k_index[2896] = 13320;
mem_k_index[2897] = 13323;
mem_k_index[2898] = 13325;
mem_k_index[2899] = 13328;
mem_k_index[2900] = 13330;
mem_k_index[2901] = 13333;
mem_k_index[2902] = 13336;
mem_k_index[2903] = 13338;
mem_k_index[2904] = 13341;
mem_k_index[2905] = 13343;
mem_k_index[2906] = 13346;
mem_k_index[2907] = 13348;
mem_k_index[2908] = 13351;
mem_k_index[2909] = 13353;
mem_k_index[2910] = 13356;
mem_k_index[2911] = 13358;
mem_k_index[2912] = 13361;
mem_k_index[2913] = 13363;
mem_k_index[2914] = 13366;
mem_k_index[2915] = 13368;
mem_k_index[2916] = 13371;
mem_k_index[2917] = 13373;
mem_k_index[2918] = 13376;
mem_k_index[2919] = 13378;
mem_k_index[2920] = 13381;
mem_k_index[2921] = 13383;
mem_k_index[2922] = 13386;
mem_k_index[2923] = 13388;
mem_k_index[2924] = 13391;
mem_k_index[2925] = 13393;
mem_k_index[2926] = 13396;
mem_k_index[2927] = 13398;
mem_k_index[2928] = 13401;
mem_k_index[2929] = 13403;
mem_k_index[2930] = 13406;
mem_k_index[2931] = 13408;
mem_k_index[2932] = 13411;
mem_k_index[2933] = 13413;
mem_k_index[2934] = 13416;
mem_k_index[2935] = 13418;
mem_k_index[2936] = 13421;
mem_k_index[2937] = 13423;
mem_k_index[2938] = 13426;
mem_k_index[2939] = 13428;
mem_k_index[2940] = 13431;
mem_k_index[2941] = 13433;
mem_k_index[2942] = 13436;
mem_k_index[2943] = 13438;
mem_k_index[2944] = 13760;
mem_k_index[2945] = 13762;
mem_k_index[2946] = 13765;
mem_k_index[2947] = 13767;
mem_k_index[2948] = 13770;
mem_k_index[2949] = 13772;
mem_k_index[2950] = 13775;
mem_k_index[2951] = 13777;
mem_k_index[2952] = 13780;
mem_k_index[2953] = 13782;
mem_k_index[2954] = 13785;
mem_k_index[2955] = 13787;
mem_k_index[2956] = 13790;
mem_k_index[2957] = 13792;
mem_k_index[2958] = 13795;
mem_k_index[2959] = 13797;
mem_k_index[2960] = 13800;
mem_k_index[2961] = 13802;
mem_k_index[2962] = 13805;
mem_k_index[2963] = 13807;
mem_k_index[2964] = 13810;
mem_k_index[2965] = 13812;
mem_k_index[2966] = 13815;
mem_k_index[2967] = 13817;
mem_k_index[2968] = 13820;
mem_k_index[2969] = 13822;
mem_k_index[2970] = 13825;
mem_k_index[2971] = 13827;
mem_k_index[2972] = 13830;
mem_k_index[2973] = 13832;
mem_k_index[2974] = 13835;
mem_k_index[2975] = 13837;
mem_k_index[2976] = 13840;
mem_k_index[2977] = 13842;
mem_k_index[2978] = 13845;
mem_k_index[2979] = 13847;
mem_k_index[2980] = 13850;
mem_k_index[2981] = 13852;
mem_k_index[2982] = 13855;
mem_k_index[2983] = 13857;
mem_k_index[2984] = 13860;
mem_k_index[2985] = 13862;
mem_k_index[2986] = 13865;
mem_k_index[2987] = 13868;
mem_k_index[2988] = 13870;
mem_k_index[2989] = 13873;
mem_k_index[2990] = 13875;
mem_k_index[2991] = 13878;
mem_k_index[2992] = 13880;
mem_k_index[2993] = 13883;
mem_k_index[2994] = 13885;
mem_k_index[2995] = 13888;
mem_k_index[2996] = 13890;
mem_k_index[2997] = 13893;
mem_k_index[2998] = 13895;
mem_k_index[2999] = 13898;
mem_k_index[3000] = 13900;
mem_k_index[3001] = 13903;
mem_k_index[3002] = 13905;
mem_k_index[3003] = 13908;
mem_k_index[3004] = 13910;
mem_k_index[3005] = 13913;
mem_k_index[3006] = 13915;
mem_k_index[3007] = 13918;
mem_k_index[3008] = 13920;
mem_k_index[3009] = 13923;
mem_k_index[3010] = 13925;
mem_k_index[3011] = 13928;
mem_k_index[3012] = 13930;
mem_k_index[3013] = 13933;
mem_k_index[3014] = 13935;
mem_k_index[3015] = 13938;
mem_k_index[3016] = 13940;
mem_k_index[3017] = 13943;
mem_k_index[3018] = 13945;
mem_k_index[3019] = 13948;
mem_k_index[3020] = 13950;
mem_k_index[3021] = 13953;
mem_k_index[3022] = 13955;
mem_k_index[3023] = 13958;
mem_k_index[3024] = 13960;
mem_k_index[3025] = 13963;
mem_k_index[3026] = 13965;
mem_k_index[3027] = 13968;
mem_k_index[3028] = 13970;
mem_k_index[3029] = 13973;
mem_k_index[3030] = 13976;
mem_k_index[3031] = 13978;
mem_k_index[3032] = 13981;
mem_k_index[3033] = 13983;
mem_k_index[3034] = 13986;
mem_k_index[3035] = 13988;
mem_k_index[3036] = 13991;
mem_k_index[3037] = 13993;
mem_k_index[3038] = 13996;
mem_k_index[3039] = 13998;
mem_k_index[3040] = 14001;
mem_k_index[3041] = 14003;
mem_k_index[3042] = 14006;
mem_k_index[3043] = 14008;
mem_k_index[3044] = 14011;
mem_k_index[3045] = 14013;
mem_k_index[3046] = 14016;
mem_k_index[3047] = 14018;
mem_k_index[3048] = 14021;
mem_k_index[3049] = 14023;
mem_k_index[3050] = 14026;
mem_k_index[3051] = 14028;
mem_k_index[3052] = 14031;
mem_k_index[3053] = 14033;
mem_k_index[3054] = 14036;
mem_k_index[3055] = 14038;
mem_k_index[3056] = 14041;
mem_k_index[3057] = 14043;
mem_k_index[3058] = 14046;
mem_k_index[3059] = 14048;
mem_k_index[3060] = 14051;
mem_k_index[3061] = 14053;
mem_k_index[3062] = 14056;
mem_k_index[3063] = 14058;
mem_k_index[3064] = 14061;
mem_k_index[3065] = 14063;
mem_k_index[3066] = 14066;
mem_k_index[3067] = 14068;
mem_k_index[3068] = 14071;
mem_k_index[3069] = 14073;
mem_k_index[3070] = 14076;
mem_k_index[3071] = 14078;
mem_k_index[3072] = 14400;
mem_k_index[3073] = 14402;
mem_k_index[3074] = 14405;
mem_k_index[3075] = 14407;
mem_k_index[3076] = 14410;
mem_k_index[3077] = 14412;
mem_k_index[3078] = 14415;
mem_k_index[3079] = 14417;
mem_k_index[3080] = 14420;
mem_k_index[3081] = 14422;
mem_k_index[3082] = 14425;
mem_k_index[3083] = 14427;
mem_k_index[3084] = 14430;
mem_k_index[3085] = 14432;
mem_k_index[3086] = 14435;
mem_k_index[3087] = 14437;
mem_k_index[3088] = 14440;
mem_k_index[3089] = 14442;
mem_k_index[3090] = 14445;
mem_k_index[3091] = 14447;
mem_k_index[3092] = 14450;
mem_k_index[3093] = 14452;
mem_k_index[3094] = 14455;
mem_k_index[3095] = 14457;
mem_k_index[3096] = 14460;
mem_k_index[3097] = 14462;
mem_k_index[3098] = 14465;
mem_k_index[3099] = 14467;
mem_k_index[3100] = 14470;
mem_k_index[3101] = 14472;
mem_k_index[3102] = 14475;
mem_k_index[3103] = 14477;
mem_k_index[3104] = 14480;
mem_k_index[3105] = 14482;
mem_k_index[3106] = 14485;
mem_k_index[3107] = 14487;
mem_k_index[3108] = 14490;
mem_k_index[3109] = 14492;
mem_k_index[3110] = 14495;
mem_k_index[3111] = 14497;
mem_k_index[3112] = 14500;
mem_k_index[3113] = 14502;
mem_k_index[3114] = 14505;
mem_k_index[3115] = 14508;
mem_k_index[3116] = 14510;
mem_k_index[3117] = 14513;
mem_k_index[3118] = 14515;
mem_k_index[3119] = 14518;
mem_k_index[3120] = 14520;
mem_k_index[3121] = 14523;
mem_k_index[3122] = 14525;
mem_k_index[3123] = 14528;
mem_k_index[3124] = 14530;
mem_k_index[3125] = 14533;
mem_k_index[3126] = 14535;
mem_k_index[3127] = 14538;
mem_k_index[3128] = 14540;
mem_k_index[3129] = 14543;
mem_k_index[3130] = 14545;
mem_k_index[3131] = 14548;
mem_k_index[3132] = 14550;
mem_k_index[3133] = 14553;
mem_k_index[3134] = 14555;
mem_k_index[3135] = 14558;
mem_k_index[3136] = 14560;
mem_k_index[3137] = 14563;
mem_k_index[3138] = 14565;
mem_k_index[3139] = 14568;
mem_k_index[3140] = 14570;
mem_k_index[3141] = 14573;
mem_k_index[3142] = 14575;
mem_k_index[3143] = 14578;
mem_k_index[3144] = 14580;
mem_k_index[3145] = 14583;
mem_k_index[3146] = 14585;
mem_k_index[3147] = 14588;
mem_k_index[3148] = 14590;
mem_k_index[3149] = 14593;
mem_k_index[3150] = 14595;
mem_k_index[3151] = 14598;
mem_k_index[3152] = 14600;
mem_k_index[3153] = 14603;
mem_k_index[3154] = 14605;
mem_k_index[3155] = 14608;
mem_k_index[3156] = 14610;
mem_k_index[3157] = 14613;
mem_k_index[3158] = 14616;
mem_k_index[3159] = 14618;
mem_k_index[3160] = 14621;
mem_k_index[3161] = 14623;
mem_k_index[3162] = 14626;
mem_k_index[3163] = 14628;
mem_k_index[3164] = 14631;
mem_k_index[3165] = 14633;
mem_k_index[3166] = 14636;
mem_k_index[3167] = 14638;
mem_k_index[3168] = 14641;
mem_k_index[3169] = 14643;
mem_k_index[3170] = 14646;
mem_k_index[3171] = 14648;
mem_k_index[3172] = 14651;
mem_k_index[3173] = 14653;
mem_k_index[3174] = 14656;
mem_k_index[3175] = 14658;
mem_k_index[3176] = 14661;
mem_k_index[3177] = 14663;
mem_k_index[3178] = 14666;
mem_k_index[3179] = 14668;
mem_k_index[3180] = 14671;
mem_k_index[3181] = 14673;
mem_k_index[3182] = 14676;
mem_k_index[3183] = 14678;
mem_k_index[3184] = 14681;
mem_k_index[3185] = 14683;
mem_k_index[3186] = 14686;
mem_k_index[3187] = 14688;
mem_k_index[3188] = 14691;
mem_k_index[3189] = 14693;
mem_k_index[3190] = 14696;
mem_k_index[3191] = 14698;
mem_k_index[3192] = 14701;
mem_k_index[3193] = 14703;
mem_k_index[3194] = 14706;
mem_k_index[3195] = 14708;
mem_k_index[3196] = 14711;
mem_k_index[3197] = 14713;
mem_k_index[3198] = 14716;
mem_k_index[3199] = 14718;
mem_k_index[3200] = 15040;
mem_k_index[3201] = 15042;
mem_k_index[3202] = 15045;
mem_k_index[3203] = 15047;
mem_k_index[3204] = 15050;
mem_k_index[3205] = 15052;
mem_k_index[3206] = 15055;
mem_k_index[3207] = 15057;
mem_k_index[3208] = 15060;
mem_k_index[3209] = 15062;
mem_k_index[3210] = 15065;
mem_k_index[3211] = 15067;
mem_k_index[3212] = 15070;
mem_k_index[3213] = 15072;
mem_k_index[3214] = 15075;
mem_k_index[3215] = 15077;
mem_k_index[3216] = 15080;
mem_k_index[3217] = 15082;
mem_k_index[3218] = 15085;
mem_k_index[3219] = 15087;
mem_k_index[3220] = 15090;
mem_k_index[3221] = 15092;
mem_k_index[3222] = 15095;
mem_k_index[3223] = 15097;
mem_k_index[3224] = 15100;
mem_k_index[3225] = 15102;
mem_k_index[3226] = 15105;
mem_k_index[3227] = 15107;
mem_k_index[3228] = 15110;
mem_k_index[3229] = 15112;
mem_k_index[3230] = 15115;
mem_k_index[3231] = 15117;
mem_k_index[3232] = 15120;
mem_k_index[3233] = 15122;
mem_k_index[3234] = 15125;
mem_k_index[3235] = 15127;
mem_k_index[3236] = 15130;
mem_k_index[3237] = 15132;
mem_k_index[3238] = 15135;
mem_k_index[3239] = 15137;
mem_k_index[3240] = 15140;
mem_k_index[3241] = 15142;
mem_k_index[3242] = 15145;
mem_k_index[3243] = 15148;
mem_k_index[3244] = 15150;
mem_k_index[3245] = 15153;
mem_k_index[3246] = 15155;
mem_k_index[3247] = 15158;
mem_k_index[3248] = 15160;
mem_k_index[3249] = 15163;
mem_k_index[3250] = 15165;
mem_k_index[3251] = 15168;
mem_k_index[3252] = 15170;
mem_k_index[3253] = 15173;
mem_k_index[3254] = 15175;
mem_k_index[3255] = 15178;
mem_k_index[3256] = 15180;
mem_k_index[3257] = 15183;
mem_k_index[3258] = 15185;
mem_k_index[3259] = 15188;
mem_k_index[3260] = 15190;
mem_k_index[3261] = 15193;
mem_k_index[3262] = 15195;
mem_k_index[3263] = 15198;
mem_k_index[3264] = 15200;
mem_k_index[3265] = 15203;
mem_k_index[3266] = 15205;
mem_k_index[3267] = 15208;
mem_k_index[3268] = 15210;
mem_k_index[3269] = 15213;
mem_k_index[3270] = 15215;
mem_k_index[3271] = 15218;
mem_k_index[3272] = 15220;
mem_k_index[3273] = 15223;
mem_k_index[3274] = 15225;
mem_k_index[3275] = 15228;
mem_k_index[3276] = 15230;
mem_k_index[3277] = 15233;
mem_k_index[3278] = 15235;
mem_k_index[3279] = 15238;
mem_k_index[3280] = 15240;
mem_k_index[3281] = 15243;
mem_k_index[3282] = 15245;
mem_k_index[3283] = 15248;
mem_k_index[3284] = 15250;
mem_k_index[3285] = 15253;
mem_k_index[3286] = 15256;
mem_k_index[3287] = 15258;
mem_k_index[3288] = 15261;
mem_k_index[3289] = 15263;
mem_k_index[3290] = 15266;
mem_k_index[3291] = 15268;
mem_k_index[3292] = 15271;
mem_k_index[3293] = 15273;
mem_k_index[3294] = 15276;
mem_k_index[3295] = 15278;
mem_k_index[3296] = 15281;
mem_k_index[3297] = 15283;
mem_k_index[3298] = 15286;
mem_k_index[3299] = 15288;
mem_k_index[3300] = 15291;
mem_k_index[3301] = 15293;
mem_k_index[3302] = 15296;
mem_k_index[3303] = 15298;
mem_k_index[3304] = 15301;
mem_k_index[3305] = 15303;
mem_k_index[3306] = 15306;
mem_k_index[3307] = 15308;
mem_k_index[3308] = 15311;
mem_k_index[3309] = 15313;
mem_k_index[3310] = 15316;
mem_k_index[3311] = 15318;
mem_k_index[3312] = 15321;
mem_k_index[3313] = 15323;
mem_k_index[3314] = 15326;
mem_k_index[3315] = 15328;
mem_k_index[3316] = 15331;
mem_k_index[3317] = 15333;
mem_k_index[3318] = 15336;
mem_k_index[3319] = 15338;
mem_k_index[3320] = 15341;
mem_k_index[3321] = 15343;
mem_k_index[3322] = 15346;
mem_k_index[3323] = 15348;
mem_k_index[3324] = 15351;
mem_k_index[3325] = 15353;
mem_k_index[3326] = 15356;
mem_k_index[3327] = 15358;
mem_k_index[3328] = 15360;
mem_k_index[3329] = 15362;
mem_k_index[3330] = 15365;
mem_k_index[3331] = 15367;
mem_k_index[3332] = 15370;
mem_k_index[3333] = 15372;
mem_k_index[3334] = 15375;
mem_k_index[3335] = 15377;
mem_k_index[3336] = 15380;
mem_k_index[3337] = 15382;
mem_k_index[3338] = 15385;
mem_k_index[3339] = 15387;
mem_k_index[3340] = 15390;
mem_k_index[3341] = 15392;
mem_k_index[3342] = 15395;
mem_k_index[3343] = 15397;
mem_k_index[3344] = 15400;
mem_k_index[3345] = 15402;
mem_k_index[3346] = 15405;
mem_k_index[3347] = 15407;
mem_k_index[3348] = 15410;
mem_k_index[3349] = 15412;
mem_k_index[3350] = 15415;
mem_k_index[3351] = 15417;
mem_k_index[3352] = 15420;
mem_k_index[3353] = 15422;
mem_k_index[3354] = 15425;
mem_k_index[3355] = 15427;
mem_k_index[3356] = 15430;
mem_k_index[3357] = 15432;
mem_k_index[3358] = 15435;
mem_k_index[3359] = 15437;
mem_k_index[3360] = 15440;
mem_k_index[3361] = 15442;
mem_k_index[3362] = 15445;
mem_k_index[3363] = 15447;
mem_k_index[3364] = 15450;
mem_k_index[3365] = 15452;
mem_k_index[3366] = 15455;
mem_k_index[3367] = 15457;
mem_k_index[3368] = 15460;
mem_k_index[3369] = 15462;
mem_k_index[3370] = 15465;
mem_k_index[3371] = 15468;
mem_k_index[3372] = 15470;
mem_k_index[3373] = 15473;
mem_k_index[3374] = 15475;
mem_k_index[3375] = 15478;
mem_k_index[3376] = 15480;
mem_k_index[3377] = 15483;
mem_k_index[3378] = 15485;
mem_k_index[3379] = 15488;
mem_k_index[3380] = 15490;
mem_k_index[3381] = 15493;
mem_k_index[3382] = 15495;
mem_k_index[3383] = 15498;
mem_k_index[3384] = 15500;
mem_k_index[3385] = 15503;
mem_k_index[3386] = 15505;
mem_k_index[3387] = 15508;
mem_k_index[3388] = 15510;
mem_k_index[3389] = 15513;
mem_k_index[3390] = 15515;
mem_k_index[3391] = 15518;
mem_k_index[3392] = 15520;
mem_k_index[3393] = 15523;
mem_k_index[3394] = 15525;
mem_k_index[3395] = 15528;
mem_k_index[3396] = 15530;
mem_k_index[3397] = 15533;
mem_k_index[3398] = 15535;
mem_k_index[3399] = 15538;
mem_k_index[3400] = 15540;
mem_k_index[3401] = 15543;
mem_k_index[3402] = 15545;
mem_k_index[3403] = 15548;
mem_k_index[3404] = 15550;
mem_k_index[3405] = 15553;
mem_k_index[3406] = 15555;
mem_k_index[3407] = 15558;
mem_k_index[3408] = 15560;
mem_k_index[3409] = 15563;
mem_k_index[3410] = 15565;
mem_k_index[3411] = 15568;
mem_k_index[3412] = 15570;
mem_k_index[3413] = 15573;
mem_k_index[3414] = 15576;
mem_k_index[3415] = 15578;
mem_k_index[3416] = 15581;
mem_k_index[3417] = 15583;
mem_k_index[3418] = 15586;
mem_k_index[3419] = 15588;
mem_k_index[3420] = 15591;
mem_k_index[3421] = 15593;
mem_k_index[3422] = 15596;
mem_k_index[3423] = 15598;
mem_k_index[3424] = 15601;
mem_k_index[3425] = 15603;
mem_k_index[3426] = 15606;
mem_k_index[3427] = 15608;
mem_k_index[3428] = 15611;
mem_k_index[3429] = 15613;
mem_k_index[3430] = 15616;
mem_k_index[3431] = 15618;
mem_k_index[3432] = 15621;
mem_k_index[3433] = 15623;
mem_k_index[3434] = 15626;
mem_k_index[3435] = 15628;
mem_k_index[3436] = 15631;
mem_k_index[3437] = 15633;
mem_k_index[3438] = 15636;
mem_k_index[3439] = 15638;
mem_k_index[3440] = 15641;
mem_k_index[3441] = 15643;
mem_k_index[3442] = 15646;
mem_k_index[3443] = 15648;
mem_k_index[3444] = 15651;
mem_k_index[3445] = 15653;
mem_k_index[3446] = 15656;
mem_k_index[3447] = 15658;
mem_k_index[3448] = 15661;
mem_k_index[3449] = 15663;
mem_k_index[3450] = 15666;
mem_k_index[3451] = 15668;
mem_k_index[3452] = 15671;
mem_k_index[3453] = 15673;
mem_k_index[3454] = 15676;
mem_k_index[3455] = 15678;
mem_k_index[3456] = 16000;
mem_k_index[3457] = 16002;
mem_k_index[3458] = 16005;
mem_k_index[3459] = 16007;
mem_k_index[3460] = 16010;
mem_k_index[3461] = 16012;
mem_k_index[3462] = 16015;
mem_k_index[3463] = 16017;
mem_k_index[3464] = 16020;
mem_k_index[3465] = 16022;
mem_k_index[3466] = 16025;
mem_k_index[3467] = 16027;
mem_k_index[3468] = 16030;
mem_k_index[3469] = 16032;
mem_k_index[3470] = 16035;
mem_k_index[3471] = 16037;
mem_k_index[3472] = 16040;
mem_k_index[3473] = 16042;
mem_k_index[3474] = 16045;
mem_k_index[3475] = 16047;
mem_k_index[3476] = 16050;
mem_k_index[3477] = 16052;
mem_k_index[3478] = 16055;
mem_k_index[3479] = 16057;
mem_k_index[3480] = 16060;
mem_k_index[3481] = 16062;
mem_k_index[3482] = 16065;
mem_k_index[3483] = 16067;
mem_k_index[3484] = 16070;
mem_k_index[3485] = 16072;
mem_k_index[3486] = 16075;
mem_k_index[3487] = 16077;
mem_k_index[3488] = 16080;
mem_k_index[3489] = 16082;
mem_k_index[3490] = 16085;
mem_k_index[3491] = 16087;
mem_k_index[3492] = 16090;
mem_k_index[3493] = 16092;
mem_k_index[3494] = 16095;
mem_k_index[3495] = 16097;
mem_k_index[3496] = 16100;
mem_k_index[3497] = 16102;
mem_k_index[3498] = 16105;
mem_k_index[3499] = 16108;
mem_k_index[3500] = 16110;
mem_k_index[3501] = 16113;
mem_k_index[3502] = 16115;
mem_k_index[3503] = 16118;
mem_k_index[3504] = 16120;
mem_k_index[3505] = 16123;
mem_k_index[3506] = 16125;
mem_k_index[3507] = 16128;
mem_k_index[3508] = 16130;
mem_k_index[3509] = 16133;
mem_k_index[3510] = 16135;
mem_k_index[3511] = 16138;
mem_k_index[3512] = 16140;
mem_k_index[3513] = 16143;
mem_k_index[3514] = 16145;
mem_k_index[3515] = 16148;
mem_k_index[3516] = 16150;
mem_k_index[3517] = 16153;
mem_k_index[3518] = 16155;
mem_k_index[3519] = 16158;
mem_k_index[3520] = 16160;
mem_k_index[3521] = 16163;
mem_k_index[3522] = 16165;
mem_k_index[3523] = 16168;
mem_k_index[3524] = 16170;
mem_k_index[3525] = 16173;
mem_k_index[3526] = 16175;
mem_k_index[3527] = 16178;
mem_k_index[3528] = 16180;
mem_k_index[3529] = 16183;
mem_k_index[3530] = 16185;
mem_k_index[3531] = 16188;
mem_k_index[3532] = 16190;
mem_k_index[3533] = 16193;
mem_k_index[3534] = 16195;
mem_k_index[3535] = 16198;
mem_k_index[3536] = 16200;
mem_k_index[3537] = 16203;
mem_k_index[3538] = 16205;
mem_k_index[3539] = 16208;
mem_k_index[3540] = 16210;
mem_k_index[3541] = 16213;
mem_k_index[3542] = 16216;
mem_k_index[3543] = 16218;
mem_k_index[3544] = 16221;
mem_k_index[3545] = 16223;
mem_k_index[3546] = 16226;
mem_k_index[3547] = 16228;
mem_k_index[3548] = 16231;
mem_k_index[3549] = 16233;
mem_k_index[3550] = 16236;
mem_k_index[3551] = 16238;
mem_k_index[3552] = 16241;
mem_k_index[3553] = 16243;
mem_k_index[3554] = 16246;
mem_k_index[3555] = 16248;
mem_k_index[3556] = 16251;
mem_k_index[3557] = 16253;
mem_k_index[3558] = 16256;
mem_k_index[3559] = 16258;
mem_k_index[3560] = 16261;
mem_k_index[3561] = 16263;
mem_k_index[3562] = 16266;
mem_k_index[3563] = 16268;
mem_k_index[3564] = 16271;
mem_k_index[3565] = 16273;
mem_k_index[3566] = 16276;
mem_k_index[3567] = 16278;
mem_k_index[3568] = 16281;
mem_k_index[3569] = 16283;
mem_k_index[3570] = 16286;
mem_k_index[3571] = 16288;
mem_k_index[3572] = 16291;
mem_k_index[3573] = 16293;
mem_k_index[3574] = 16296;
mem_k_index[3575] = 16298;
mem_k_index[3576] = 16301;
mem_k_index[3577] = 16303;
mem_k_index[3578] = 16306;
mem_k_index[3579] = 16308;
mem_k_index[3580] = 16311;
mem_k_index[3581] = 16313;
mem_k_index[3582] = 16316;
mem_k_index[3583] = 16318;
mem_k_index[3584] = 16640;
mem_k_index[3585] = 16642;
mem_k_index[3586] = 16645;
mem_k_index[3587] = 16647;
mem_k_index[3588] = 16650;
mem_k_index[3589] = 16652;
mem_k_index[3590] = 16655;
mem_k_index[3591] = 16657;
mem_k_index[3592] = 16660;
mem_k_index[3593] = 16662;
mem_k_index[3594] = 16665;
mem_k_index[3595] = 16667;
mem_k_index[3596] = 16670;
mem_k_index[3597] = 16672;
mem_k_index[3598] = 16675;
mem_k_index[3599] = 16677;
mem_k_index[3600] = 16680;
mem_k_index[3601] = 16682;
mem_k_index[3602] = 16685;
mem_k_index[3603] = 16687;
mem_k_index[3604] = 16690;
mem_k_index[3605] = 16692;
mem_k_index[3606] = 16695;
mem_k_index[3607] = 16697;
mem_k_index[3608] = 16700;
mem_k_index[3609] = 16702;
mem_k_index[3610] = 16705;
mem_k_index[3611] = 16707;
mem_k_index[3612] = 16710;
mem_k_index[3613] = 16712;
mem_k_index[3614] = 16715;
mem_k_index[3615] = 16717;
mem_k_index[3616] = 16720;
mem_k_index[3617] = 16722;
mem_k_index[3618] = 16725;
mem_k_index[3619] = 16727;
mem_k_index[3620] = 16730;
mem_k_index[3621] = 16732;
mem_k_index[3622] = 16735;
mem_k_index[3623] = 16737;
mem_k_index[3624] = 16740;
mem_k_index[3625] = 16742;
mem_k_index[3626] = 16745;
mem_k_index[3627] = 16748;
mem_k_index[3628] = 16750;
mem_k_index[3629] = 16753;
mem_k_index[3630] = 16755;
mem_k_index[3631] = 16758;
mem_k_index[3632] = 16760;
mem_k_index[3633] = 16763;
mem_k_index[3634] = 16765;
mem_k_index[3635] = 16768;
mem_k_index[3636] = 16770;
mem_k_index[3637] = 16773;
mem_k_index[3638] = 16775;
mem_k_index[3639] = 16778;
mem_k_index[3640] = 16780;
mem_k_index[3641] = 16783;
mem_k_index[3642] = 16785;
mem_k_index[3643] = 16788;
mem_k_index[3644] = 16790;
mem_k_index[3645] = 16793;
mem_k_index[3646] = 16795;
mem_k_index[3647] = 16798;
mem_k_index[3648] = 16800;
mem_k_index[3649] = 16803;
mem_k_index[3650] = 16805;
mem_k_index[3651] = 16808;
mem_k_index[3652] = 16810;
mem_k_index[3653] = 16813;
mem_k_index[3654] = 16815;
mem_k_index[3655] = 16818;
mem_k_index[3656] = 16820;
mem_k_index[3657] = 16823;
mem_k_index[3658] = 16825;
mem_k_index[3659] = 16828;
mem_k_index[3660] = 16830;
mem_k_index[3661] = 16833;
mem_k_index[3662] = 16835;
mem_k_index[3663] = 16838;
mem_k_index[3664] = 16840;
mem_k_index[3665] = 16843;
mem_k_index[3666] = 16845;
mem_k_index[3667] = 16848;
mem_k_index[3668] = 16850;
mem_k_index[3669] = 16853;
mem_k_index[3670] = 16856;
mem_k_index[3671] = 16858;
mem_k_index[3672] = 16861;
mem_k_index[3673] = 16863;
mem_k_index[3674] = 16866;
mem_k_index[3675] = 16868;
mem_k_index[3676] = 16871;
mem_k_index[3677] = 16873;
mem_k_index[3678] = 16876;
mem_k_index[3679] = 16878;
mem_k_index[3680] = 16881;
mem_k_index[3681] = 16883;
mem_k_index[3682] = 16886;
mem_k_index[3683] = 16888;
mem_k_index[3684] = 16891;
mem_k_index[3685] = 16893;
mem_k_index[3686] = 16896;
mem_k_index[3687] = 16898;
mem_k_index[3688] = 16901;
mem_k_index[3689] = 16903;
mem_k_index[3690] = 16906;
mem_k_index[3691] = 16908;
mem_k_index[3692] = 16911;
mem_k_index[3693] = 16913;
mem_k_index[3694] = 16916;
mem_k_index[3695] = 16918;
mem_k_index[3696] = 16921;
mem_k_index[3697] = 16923;
mem_k_index[3698] = 16926;
mem_k_index[3699] = 16928;
mem_k_index[3700] = 16931;
mem_k_index[3701] = 16933;
mem_k_index[3702] = 16936;
mem_k_index[3703] = 16938;
mem_k_index[3704] = 16941;
mem_k_index[3705] = 16943;
mem_k_index[3706] = 16946;
mem_k_index[3707] = 16948;
mem_k_index[3708] = 16951;
mem_k_index[3709] = 16953;
mem_k_index[3710] = 16956;
mem_k_index[3711] = 16958;
mem_k_index[3712] = 17280;
mem_k_index[3713] = 17282;
mem_k_index[3714] = 17285;
mem_k_index[3715] = 17287;
mem_k_index[3716] = 17290;
mem_k_index[3717] = 17292;
mem_k_index[3718] = 17295;
mem_k_index[3719] = 17297;
mem_k_index[3720] = 17300;
mem_k_index[3721] = 17302;
mem_k_index[3722] = 17305;
mem_k_index[3723] = 17307;
mem_k_index[3724] = 17310;
mem_k_index[3725] = 17312;
mem_k_index[3726] = 17315;
mem_k_index[3727] = 17317;
mem_k_index[3728] = 17320;
mem_k_index[3729] = 17322;
mem_k_index[3730] = 17325;
mem_k_index[3731] = 17327;
mem_k_index[3732] = 17330;
mem_k_index[3733] = 17332;
mem_k_index[3734] = 17335;
mem_k_index[3735] = 17337;
mem_k_index[3736] = 17340;
mem_k_index[3737] = 17342;
mem_k_index[3738] = 17345;
mem_k_index[3739] = 17347;
mem_k_index[3740] = 17350;
mem_k_index[3741] = 17352;
mem_k_index[3742] = 17355;
mem_k_index[3743] = 17357;
mem_k_index[3744] = 17360;
mem_k_index[3745] = 17362;
mem_k_index[3746] = 17365;
mem_k_index[3747] = 17367;
mem_k_index[3748] = 17370;
mem_k_index[3749] = 17372;
mem_k_index[3750] = 17375;
mem_k_index[3751] = 17377;
mem_k_index[3752] = 17380;
mem_k_index[3753] = 17382;
mem_k_index[3754] = 17385;
mem_k_index[3755] = 17388;
mem_k_index[3756] = 17390;
mem_k_index[3757] = 17393;
mem_k_index[3758] = 17395;
mem_k_index[3759] = 17398;
mem_k_index[3760] = 17400;
mem_k_index[3761] = 17403;
mem_k_index[3762] = 17405;
mem_k_index[3763] = 17408;
mem_k_index[3764] = 17410;
mem_k_index[3765] = 17413;
mem_k_index[3766] = 17415;
mem_k_index[3767] = 17418;
mem_k_index[3768] = 17420;
mem_k_index[3769] = 17423;
mem_k_index[3770] = 17425;
mem_k_index[3771] = 17428;
mem_k_index[3772] = 17430;
mem_k_index[3773] = 17433;
mem_k_index[3774] = 17435;
mem_k_index[3775] = 17438;
mem_k_index[3776] = 17440;
mem_k_index[3777] = 17443;
mem_k_index[3778] = 17445;
mem_k_index[3779] = 17448;
mem_k_index[3780] = 17450;
mem_k_index[3781] = 17453;
mem_k_index[3782] = 17455;
mem_k_index[3783] = 17458;
mem_k_index[3784] = 17460;
mem_k_index[3785] = 17463;
mem_k_index[3786] = 17465;
mem_k_index[3787] = 17468;
mem_k_index[3788] = 17470;
mem_k_index[3789] = 17473;
mem_k_index[3790] = 17475;
mem_k_index[3791] = 17478;
mem_k_index[3792] = 17480;
mem_k_index[3793] = 17483;
mem_k_index[3794] = 17485;
mem_k_index[3795] = 17488;
mem_k_index[3796] = 17490;
mem_k_index[3797] = 17493;
mem_k_index[3798] = 17496;
mem_k_index[3799] = 17498;
mem_k_index[3800] = 17501;
mem_k_index[3801] = 17503;
mem_k_index[3802] = 17506;
mem_k_index[3803] = 17508;
mem_k_index[3804] = 17511;
mem_k_index[3805] = 17513;
mem_k_index[3806] = 17516;
mem_k_index[3807] = 17518;
mem_k_index[3808] = 17521;
mem_k_index[3809] = 17523;
mem_k_index[3810] = 17526;
mem_k_index[3811] = 17528;
mem_k_index[3812] = 17531;
mem_k_index[3813] = 17533;
mem_k_index[3814] = 17536;
mem_k_index[3815] = 17538;
mem_k_index[3816] = 17541;
mem_k_index[3817] = 17543;
mem_k_index[3818] = 17546;
mem_k_index[3819] = 17548;
mem_k_index[3820] = 17551;
mem_k_index[3821] = 17553;
mem_k_index[3822] = 17556;
mem_k_index[3823] = 17558;
mem_k_index[3824] = 17561;
mem_k_index[3825] = 17563;
mem_k_index[3826] = 17566;
mem_k_index[3827] = 17568;
mem_k_index[3828] = 17571;
mem_k_index[3829] = 17573;
mem_k_index[3830] = 17576;
mem_k_index[3831] = 17578;
mem_k_index[3832] = 17581;
mem_k_index[3833] = 17583;
mem_k_index[3834] = 17586;
mem_k_index[3835] = 17588;
mem_k_index[3836] = 17591;
mem_k_index[3837] = 17593;
mem_k_index[3838] = 17596;
mem_k_index[3839] = 17598;
mem_k_index[3840] = 17920;
mem_k_index[3841] = 17922;
mem_k_index[3842] = 17925;
mem_k_index[3843] = 17927;
mem_k_index[3844] = 17930;
mem_k_index[3845] = 17932;
mem_k_index[3846] = 17935;
mem_k_index[3847] = 17937;
mem_k_index[3848] = 17940;
mem_k_index[3849] = 17942;
mem_k_index[3850] = 17945;
mem_k_index[3851] = 17947;
mem_k_index[3852] = 17950;
mem_k_index[3853] = 17952;
mem_k_index[3854] = 17955;
mem_k_index[3855] = 17957;
mem_k_index[3856] = 17960;
mem_k_index[3857] = 17962;
mem_k_index[3858] = 17965;
mem_k_index[3859] = 17967;
mem_k_index[3860] = 17970;
mem_k_index[3861] = 17972;
mem_k_index[3862] = 17975;
mem_k_index[3863] = 17977;
mem_k_index[3864] = 17980;
mem_k_index[3865] = 17982;
mem_k_index[3866] = 17985;
mem_k_index[3867] = 17987;
mem_k_index[3868] = 17990;
mem_k_index[3869] = 17992;
mem_k_index[3870] = 17995;
mem_k_index[3871] = 17997;
mem_k_index[3872] = 18000;
mem_k_index[3873] = 18002;
mem_k_index[3874] = 18005;
mem_k_index[3875] = 18007;
mem_k_index[3876] = 18010;
mem_k_index[3877] = 18012;
mem_k_index[3878] = 18015;
mem_k_index[3879] = 18017;
mem_k_index[3880] = 18020;
mem_k_index[3881] = 18022;
mem_k_index[3882] = 18025;
mem_k_index[3883] = 18028;
mem_k_index[3884] = 18030;
mem_k_index[3885] = 18033;
mem_k_index[3886] = 18035;
mem_k_index[3887] = 18038;
mem_k_index[3888] = 18040;
mem_k_index[3889] = 18043;
mem_k_index[3890] = 18045;
mem_k_index[3891] = 18048;
mem_k_index[3892] = 18050;
mem_k_index[3893] = 18053;
mem_k_index[3894] = 18055;
mem_k_index[3895] = 18058;
mem_k_index[3896] = 18060;
mem_k_index[3897] = 18063;
mem_k_index[3898] = 18065;
mem_k_index[3899] = 18068;
mem_k_index[3900] = 18070;
mem_k_index[3901] = 18073;
mem_k_index[3902] = 18075;
mem_k_index[3903] = 18078;
mem_k_index[3904] = 18080;
mem_k_index[3905] = 18083;
mem_k_index[3906] = 18085;
mem_k_index[3907] = 18088;
mem_k_index[3908] = 18090;
mem_k_index[3909] = 18093;
mem_k_index[3910] = 18095;
mem_k_index[3911] = 18098;
mem_k_index[3912] = 18100;
mem_k_index[3913] = 18103;
mem_k_index[3914] = 18105;
mem_k_index[3915] = 18108;
mem_k_index[3916] = 18110;
mem_k_index[3917] = 18113;
mem_k_index[3918] = 18115;
mem_k_index[3919] = 18118;
mem_k_index[3920] = 18120;
mem_k_index[3921] = 18123;
mem_k_index[3922] = 18125;
mem_k_index[3923] = 18128;
mem_k_index[3924] = 18130;
mem_k_index[3925] = 18133;
mem_k_index[3926] = 18136;
mem_k_index[3927] = 18138;
mem_k_index[3928] = 18141;
mem_k_index[3929] = 18143;
mem_k_index[3930] = 18146;
mem_k_index[3931] = 18148;
mem_k_index[3932] = 18151;
mem_k_index[3933] = 18153;
mem_k_index[3934] = 18156;
mem_k_index[3935] = 18158;
mem_k_index[3936] = 18161;
mem_k_index[3937] = 18163;
mem_k_index[3938] = 18166;
mem_k_index[3939] = 18168;
mem_k_index[3940] = 18171;
mem_k_index[3941] = 18173;
mem_k_index[3942] = 18176;
mem_k_index[3943] = 18178;
mem_k_index[3944] = 18181;
mem_k_index[3945] = 18183;
mem_k_index[3946] = 18186;
mem_k_index[3947] = 18188;
mem_k_index[3948] = 18191;
mem_k_index[3949] = 18193;
mem_k_index[3950] = 18196;
mem_k_index[3951] = 18198;
mem_k_index[3952] = 18201;
mem_k_index[3953] = 18203;
mem_k_index[3954] = 18206;
mem_k_index[3955] = 18208;
mem_k_index[3956] = 18211;
mem_k_index[3957] = 18213;
mem_k_index[3958] = 18216;
mem_k_index[3959] = 18218;
mem_k_index[3960] = 18221;
mem_k_index[3961] = 18223;
mem_k_index[3962] = 18226;
mem_k_index[3963] = 18228;
mem_k_index[3964] = 18231;
mem_k_index[3965] = 18233;
mem_k_index[3966] = 18236;
mem_k_index[3967] = 18238;
mem_k_index[3968] = 18560;
mem_k_index[3969] = 18562;
mem_k_index[3970] = 18565;
mem_k_index[3971] = 18567;
mem_k_index[3972] = 18570;
mem_k_index[3973] = 18572;
mem_k_index[3974] = 18575;
mem_k_index[3975] = 18577;
mem_k_index[3976] = 18580;
mem_k_index[3977] = 18582;
mem_k_index[3978] = 18585;
mem_k_index[3979] = 18587;
mem_k_index[3980] = 18590;
mem_k_index[3981] = 18592;
mem_k_index[3982] = 18595;
mem_k_index[3983] = 18597;
mem_k_index[3984] = 18600;
mem_k_index[3985] = 18602;
mem_k_index[3986] = 18605;
mem_k_index[3987] = 18607;
mem_k_index[3988] = 18610;
mem_k_index[3989] = 18612;
mem_k_index[3990] = 18615;
mem_k_index[3991] = 18617;
mem_k_index[3992] = 18620;
mem_k_index[3993] = 18622;
mem_k_index[3994] = 18625;
mem_k_index[3995] = 18627;
mem_k_index[3996] = 18630;
mem_k_index[3997] = 18632;
mem_k_index[3998] = 18635;
mem_k_index[3999] = 18637;
mem_k_index[4000] = 18640;
mem_k_index[4001] = 18642;
mem_k_index[4002] = 18645;
mem_k_index[4003] = 18647;
mem_k_index[4004] = 18650;
mem_k_index[4005] = 18652;
mem_k_index[4006] = 18655;
mem_k_index[4007] = 18657;
mem_k_index[4008] = 18660;
mem_k_index[4009] = 18662;
mem_k_index[4010] = 18665;
mem_k_index[4011] = 18668;
mem_k_index[4012] = 18670;
mem_k_index[4013] = 18673;
mem_k_index[4014] = 18675;
mem_k_index[4015] = 18678;
mem_k_index[4016] = 18680;
mem_k_index[4017] = 18683;
mem_k_index[4018] = 18685;
mem_k_index[4019] = 18688;
mem_k_index[4020] = 18690;
mem_k_index[4021] = 18693;
mem_k_index[4022] = 18695;
mem_k_index[4023] = 18698;
mem_k_index[4024] = 18700;
mem_k_index[4025] = 18703;
mem_k_index[4026] = 18705;
mem_k_index[4027] = 18708;
mem_k_index[4028] = 18710;
mem_k_index[4029] = 18713;
mem_k_index[4030] = 18715;
mem_k_index[4031] = 18718;
mem_k_index[4032] = 18720;
mem_k_index[4033] = 18723;
mem_k_index[4034] = 18725;
mem_k_index[4035] = 18728;
mem_k_index[4036] = 18730;
mem_k_index[4037] = 18733;
mem_k_index[4038] = 18735;
mem_k_index[4039] = 18738;
mem_k_index[4040] = 18740;
mem_k_index[4041] = 18743;
mem_k_index[4042] = 18745;
mem_k_index[4043] = 18748;
mem_k_index[4044] = 18750;
mem_k_index[4045] = 18753;
mem_k_index[4046] = 18755;
mem_k_index[4047] = 18758;
mem_k_index[4048] = 18760;
mem_k_index[4049] = 18763;
mem_k_index[4050] = 18765;
mem_k_index[4051] = 18768;
mem_k_index[4052] = 18770;
mem_k_index[4053] = 18773;
mem_k_index[4054] = 18776;
mem_k_index[4055] = 18778;
mem_k_index[4056] = 18781;
mem_k_index[4057] = 18783;
mem_k_index[4058] = 18786;
mem_k_index[4059] = 18788;
mem_k_index[4060] = 18791;
mem_k_index[4061] = 18793;
mem_k_index[4062] = 18796;
mem_k_index[4063] = 18798;
mem_k_index[4064] = 18801;
mem_k_index[4065] = 18803;
mem_k_index[4066] = 18806;
mem_k_index[4067] = 18808;
mem_k_index[4068] = 18811;
mem_k_index[4069] = 18813;
mem_k_index[4070] = 18816;
mem_k_index[4071] = 18818;
mem_k_index[4072] = 18821;
mem_k_index[4073] = 18823;
mem_k_index[4074] = 18826;
mem_k_index[4075] = 18828;
mem_k_index[4076] = 18831;
mem_k_index[4077] = 18833;
mem_k_index[4078] = 18836;
mem_k_index[4079] = 18838;
mem_k_index[4080] = 18841;
mem_k_index[4081] = 18843;
mem_k_index[4082] = 18846;
mem_k_index[4083] = 18848;
mem_k_index[4084] = 18851;
mem_k_index[4085] = 18853;
mem_k_index[4086] = 18856;
mem_k_index[4087] = 18858;
mem_k_index[4088] = 18861;
mem_k_index[4089] = 18863;
mem_k_index[4090] = 18866;
mem_k_index[4091] = 18868;
mem_k_index[4092] = 18871;
mem_k_index[4093] = 18873;
mem_k_index[4094] = 18876;
mem_k_index[4095] = 18878;
mem_k_index[4096] = 19200;
mem_k_index[4097] = 19202;
mem_k_index[4098] = 19205;
mem_k_index[4099] = 19207;
mem_k_index[4100] = 19210;
mem_k_index[4101] = 19212;
mem_k_index[4102] = 19215;
mem_k_index[4103] = 19217;
mem_k_index[4104] = 19220;
mem_k_index[4105] = 19222;
mem_k_index[4106] = 19225;
mem_k_index[4107] = 19227;
mem_k_index[4108] = 19230;
mem_k_index[4109] = 19232;
mem_k_index[4110] = 19235;
mem_k_index[4111] = 19237;
mem_k_index[4112] = 19240;
mem_k_index[4113] = 19242;
mem_k_index[4114] = 19245;
mem_k_index[4115] = 19247;
mem_k_index[4116] = 19250;
mem_k_index[4117] = 19252;
mem_k_index[4118] = 19255;
mem_k_index[4119] = 19257;
mem_k_index[4120] = 19260;
mem_k_index[4121] = 19262;
mem_k_index[4122] = 19265;
mem_k_index[4123] = 19267;
mem_k_index[4124] = 19270;
mem_k_index[4125] = 19272;
mem_k_index[4126] = 19275;
mem_k_index[4127] = 19277;
mem_k_index[4128] = 19280;
mem_k_index[4129] = 19282;
mem_k_index[4130] = 19285;
mem_k_index[4131] = 19287;
mem_k_index[4132] = 19290;
mem_k_index[4133] = 19292;
mem_k_index[4134] = 19295;
mem_k_index[4135] = 19297;
mem_k_index[4136] = 19300;
mem_k_index[4137] = 19302;
mem_k_index[4138] = 19305;
mem_k_index[4139] = 19308;
mem_k_index[4140] = 19310;
mem_k_index[4141] = 19313;
mem_k_index[4142] = 19315;
mem_k_index[4143] = 19318;
mem_k_index[4144] = 19320;
mem_k_index[4145] = 19323;
mem_k_index[4146] = 19325;
mem_k_index[4147] = 19328;
mem_k_index[4148] = 19330;
mem_k_index[4149] = 19333;
mem_k_index[4150] = 19335;
mem_k_index[4151] = 19338;
mem_k_index[4152] = 19340;
mem_k_index[4153] = 19343;
mem_k_index[4154] = 19345;
mem_k_index[4155] = 19348;
mem_k_index[4156] = 19350;
mem_k_index[4157] = 19353;
mem_k_index[4158] = 19355;
mem_k_index[4159] = 19358;
mem_k_index[4160] = 19360;
mem_k_index[4161] = 19363;
mem_k_index[4162] = 19365;
mem_k_index[4163] = 19368;
mem_k_index[4164] = 19370;
mem_k_index[4165] = 19373;
mem_k_index[4166] = 19375;
mem_k_index[4167] = 19378;
mem_k_index[4168] = 19380;
mem_k_index[4169] = 19383;
mem_k_index[4170] = 19385;
mem_k_index[4171] = 19388;
mem_k_index[4172] = 19390;
mem_k_index[4173] = 19393;
mem_k_index[4174] = 19395;
mem_k_index[4175] = 19398;
mem_k_index[4176] = 19400;
mem_k_index[4177] = 19403;
mem_k_index[4178] = 19405;
mem_k_index[4179] = 19408;
mem_k_index[4180] = 19410;
mem_k_index[4181] = 19413;
mem_k_index[4182] = 19416;
mem_k_index[4183] = 19418;
mem_k_index[4184] = 19421;
mem_k_index[4185] = 19423;
mem_k_index[4186] = 19426;
mem_k_index[4187] = 19428;
mem_k_index[4188] = 19431;
mem_k_index[4189] = 19433;
mem_k_index[4190] = 19436;
mem_k_index[4191] = 19438;
mem_k_index[4192] = 19441;
mem_k_index[4193] = 19443;
mem_k_index[4194] = 19446;
mem_k_index[4195] = 19448;
mem_k_index[4196] = 19451;
mem_k_index[4197] = 19453;
mem_k_index[4198] = 19456;
mem_k_index[4199] = 19458;
mem_k_index[4200] = 19461;
mem_k_index[4201] = 19463;
mem_k_index[4202] = 19466;
mem_k_index[4203] = 19468;
mem_k_index[4204] = 19471;
mem_k_index[4205] = 19473;
mem_k_index[4206] = 19476;
mem_k_index[4207] = 19478;
mem_k_index[4208] = 19481;
mem_k_index[4209] = 19483;
mem_k_index[4210] = 19486;
mem_k_index[4211] = 19488;
mem_k_index[4212] = 19491;
mem_k_index[4213] = 19493;
mem_k_index[4214] = 19496;
mem_k_index[4215] = 19498;
mem_k_index[4216] = 19501;
mem_k_index[4217] = 19503;
mem_k_index[4218] = 19506;
mem_k_index[4219] = 19508;
mem_k_index[4220] = 19511;
mem_k_index[4221] = 19513;
mem_k_index[4222] = 19516;
mem_k_index[4223] = 19518;
mem_k_index[4224] = 19840;
mem_k_index[4225] = 19842;
mem_k_index[4226] = 19845;
mem_k_index[4227] = 19847;
mem_k_index[4228] = 19850;
mem_k_index[4229] = 19852;
mem_k_index[4230] = 19855;
mem_k_index[4231] = 19857;
mem_k_index[4232] = 19860;
mem_k_index[4233] = 19862;
mem_k_index[4234] = 19865;
mem_k_index[4235] = 19867;
mem_k_index[4236] = 19870;
mem_k_index[4237] = 19872;
mem_k_index[4238] = 19875;
mem_k_index[4239] = 19877;
mem_k_index[4240] = 19880;
mem_k_index[4241] = 19882;
mem_k_index[4242] = 19885;
mem_k_index[4243] = 19887;
mem_k_index[4244] = 19890;
mem_k_index[4245] = 19892;
mem_k_index[4246] = 19895;
mem_k_index[4247] = 19897;
mem_k_index[4248] = 19900;
mem_k_index[4249] = 19902;
mem_k_index[4250] = 19905;
mem_k_index[4251] = 19907;
mem_k_index[4252] = 19910;
mem_k_index[4253] = 19912;
mem_k_index[4254] = 19915;
mem_k_index[4255] = 19917;
mem_k_index[4256] = 19920;
mem_k_index[4257] = 19922;
mem_k_index[4258] = 19925;
mem_k_index[4259] = 19927;
mem_k_index[4260] = 19930;
mem_k_index[4261] = 19932;
mem_k_index[4262] = 19935;
mem_k_index[4263] = 19937;
mem_k_index[4264] = 19940;
mem_k_index[4265] = 19942;
mem_k_index[4266] = 19945;
mem_k_index[4267] = 19948;
mem_k_index[4268] = 19950;
mem_k_index[4269] = 19953;
mem_k_index[4270] = 19955;
mem_k_index[4271] = 19958;
mem_k_index[4272] = 19960;
mem_k_index[4273] = 19963;
mem_k_index[4274] = 19965;
mem_k_index[4275] = 19968;
mem_k_index[4276] = 19970;
mem_k_index[4277] = 19973;
mem_k_index[4278] = 19975;
mem_k_index[4279] = 19978;
mem_k_index[4280] = 19980;
mem_k_index[4281] = 19983;
mem_k_index[4282] = 19985;
mem_k_index[4283] = 19988;
mem_k_index[4284] = 19990;
mem_k_index[4285] = 19993;
mem_k_index[4286] = 19995;
mem_k_index[4287] = 19998;
mem_k_index[4288] = 20000;
mem_k_index[4289] = 20003;
mem_k_index[4290] = 20005;
mem_k_index[4291] = 20008;
mem_k_index[4292] = 20010;
mem_k_index[4293] = 20013;
mem_k_index[4294] = 20015;
mem_k_index[4295] = 20018;
mem_k_index[4296] = 20020;
mem_k_index[4297] = 20023;
mem_k_index[4298] = 20025;
mem_k_index[4299] = 20028;
mem_k_index[4300] = 20030;
mem_k_index[4301] = 20033;
mem_k_index[4302] = 20035;
mem_k_index[4303] = 20038;
mem_k_index[4304] = 20040;
mem_k_index[4305] = 20043;
mem_k_index[4306] = 20045;
mem_k_index[4307] = 20048;
mem_k_index[4308] = 20050;
mem_k_index[4309] = 20053;
mem_k_index[4310] = 20056;
mem_k_index[4311] = 20058;
mem_k_index[4312] = 20061;
mem_k_index[4313] = 20063;
mem_k_index[4314] = 20066;
mem_k_index[4315] = 20068;
mem_k_index[4316] = 20071;
mem_k_index[4317] = 20073;
mem_k_index[4318] = 20076;
mem_k_index[4319] = 20078;
mem_k_index[4320] = 20081;
mem_k_index[4321] = 20083;
mem_k_index[4322] = 20086;
mem_k_index[4323] = 20088;
mem_k_index[4324] = 20091;
mem_k_index[4325] = 20093;
mem_k_index[4326] = 20096;
mem_k_index[4327] = 20098;
mem_k_index[4328] = 20101;
mem_k_index[4329] = 20103;
mem_k_index[4330] = 20106;
mem_k_index[4331] = 20108;
mem_k_index[4332] = 20111;
mem_k_index[4333] = 20113;
mem_k_index[4334] = 20116;
mem_k_index[4335] = 20118;
mem_k_index[4336] = 20121;
mem_k_index[4337] = 20123;
mem_k_index[4338] = 20126;
mem_k_index[4339] = 20128;
mem_k_index[4340] = 20131;
mem_k_index[4341] = 20133;
mem_k_index[4342] = 20136;
mem_k_index[4343] = 20138;
mem_k_index[4344] = 20141;
mem_k_index[4345] = 20143;
mem_k_index[4346] = 20146;
mem_k_index[4347] = 20148;
mem_k_index[4348] = 20151;
mem_k_index[4349] = 20153;
mem_k_index[4350] = 20156;
mem_k_index[4351] = 20158;
mem_k_index[4352] = 20160;
mem_k_index[4353] = 20162;
mem_k_index[4354] = 20165;
mem_k_index[4355] = 20167;
mem_k_index[4356] = 20170;
mem_k_index[4357] = 20172;
mem_k_index[4358] = 20175;
mem_k_index[4359] = 20177;
mem_k_index[4360] = 20180;
mem_k_index[4361] = 20182;
mem_k_index[4362] = 20185;
mem_k_index[4363] = 20187;
mem_k_index[4364] = 20190;
mem_k_index[4365] = 20192;
mem_k_index[4366] = 20195;
mem_k_index[4367] = 20197;
mem_k_index[4368] = 20200;
mem_k_index[4369] = 20202;
mem_k_index[4370] = 20205;
mem_k_index[4371] = 20207;
mem_k_index[4372] = 20210;
mem_k_index[4373] = 20212;
mem_k_index[4374] = 20215;
mem_k_index[4375] = 20217;
mem_k_index[4376] = 20220;
mem_k_index[4377] = 20222;
mem_k_index[4378] = 20225;
mem_k_index[4379] = 20227;
mem_k_index[4380] = 20230;
mem_k_index[4381] = 20232;
mem_k_index[4382] = 20235;
mem_k_index[4383] = 20237;
mem_k_index[4384] = 20240;
mem_k_index[4385] = 20242;
mem_k_index[4386] = 20245;
mem_k_index[4387] = 20247;
mem_k_index[4388] = 20250;
mem_k_index[4389] = 20252;
mem_k_index[4390] = 20255;
mem_k_index[4391] = 20257;
mem_k_index[4392] = 20260;
mem_k_index[4393] = 20262;
mem_k_index[4394] = 20265;
mem_k_index[4395] = 20268;
mem_k_index[4396] = 20270;
mem_k_index[4397] = 20273;
mem_k_index[4398] = 20275;
mem_k_index[4399] = 20278;
mem_k_index[4400] = 20280;
mem_k_index[4401] = 20283;
mem_k_index[4402] = 20285;
mem_k_index[4403] = 20288;
mem_k_index[4404] = 20290;
mem_k_index[4405] = 20293;
mem_k_index[4406] = 20295;
mem_k_index[4407] = 20298;
mem_k_index[4408] = 20300;
mem_k_index[4409] = 20303;
mem_k_index[4410] = 20305;
mem_k_index[4411] = 20308;
mem_k_index[4412] = 20310;
mem_k_index[4413] = 20313;
mem_k_index[4414] = 20315;
mem_k_index[4415] = 20318;
mem_k_index[4416] = 20320;
mem_k_index[4417] = 20323;
mem_k_index[4418] = 20325;
mem_k_index[4419] = 20328;
mem_k_index[4420] = 20330;
mem_k_index[4421] = 20333;
mem_k_index[4422] = 20335;
mem_k_index[4423] = 20338;
mem_k_index[4424] = 20340;
mem_k_index[4425] = 20343;
mem_k_index[4426] = 20345;
mem_k_index[4427] = 20348;
mem_k_index[4428] = 20350;
mem_k_index[4429] = 20353;
mem_k_index[4430] = 20355;
mem_k_index[4431] = 20358;
mem_k_index[4432] = 20360;
mem_k_index[4433] = 20363;
mem_k_index[4434] = 20365;
mem_k_index[4435] = 20368;
mem_k_index[4436] = 20370;
mem_k_index[4437] = 20373;
mem_k_index[4438] = 20376;
mem_k_index[4439] = 20378;
mem_k_index[4440] = 20381;
mem_k_index[4441] = 20383;
mem_k_index[4442] = 20386;
mem_k_index[4443] = 20388;
mem_k_index[4444] = 20391;
mem_k_index[4445] = 20393;
mem_k_index[4446] = 20396;
mem_k_index[4447] = 20398;
mem_k_index[4448] = 20401;
mem_k_index[4449] = 20403;
mem_k_index[4450] = 20406;
mem_k_index[4451] = 20408;
mem_k_index[4452] = 20411;
mem_k_index[4453] = 20413;
mem_k_index[4454] = 20416;
mem_k_index[4455] = 20418;
mem_k_index[4456] = 20421;
mem_k_index[4457] = 20423;
mem_k_index[4458] = 20426;
mem_k_index[4459] = 20428;
mem_k_index[4460] = 20431;
mem_k_index[4461] = 20433;
mem_k_index[4462] = 20436;
mem_k_index[4463] = 20438;
mem_k_index[4464] = 20441;
mem_k_index[4465] = 20443;
mem_k_index[4466] = 20446;
mem_k_index[4467] = 20448;
mem_k_index[4468] = 20451;
mem_k_index[4469] = 20453;
mem_k_index[4470] = 20456;
mem_k_index[4471] = 20458;
mem_k_index[4472] = 20461;
mem_k_index[4473] = 20463;
mem_k_index[4474] = 20466;
mem_k_index[4475] = 20468;
mem_k_index[4476] = 20471;
mem_k_index[4477] = 20473;
mem_k_index[4478] = 20476;
mem_k_index[4479] = 20478;
mem_k_index[4480] = 20800;
mem_k_index[4481] = 20802;
mem_k_index[4482] = 20805;
mem_k_index[4483] = 20807;
mem_k_index[4484] = 20810;
mem_k_index[4485] = 20812;
mem_k_index[4486] = 20815;
mem_k_index[4487] = 20817;
mem_k_index[4488] = 20820;
mem_k_index[4489] = 20822;
mem_k_index[4490] = 20825;
mem_k_index[4491] = 20827;
mem_k_index[4492] = 20830;
mem_k_index[4493] = 20832;
mem_k_index[4494] = 20835;
mem_k_index[4495] = 20837;
mem_k_index[4496] = 20840;
mem_k_index[4497] = 20842;
mem_k_index[4498] = 20845;
mem_k_index[4499] = 20847;
mem_k_index[4500] = 20850;
mem_k_index[4501] = 20852;
mem_k_index[4502] = 20855;
mem_k_index[4503] = 20857;
mem_k_index[4504] = 20860;
mem_k_index[4505] = 20862;
mem_k_index[4506] = 20865;
mem_k_index[4507] = 20867;
mem_k_index[4508] = 20870;
mem_k_index[4509] = 20872;
mem_k_index[4510] = 20875;
mem_k_index[4511] = 20877;
mem_k_index[4512] = 20880;
mem_k_index[4513] = 20882;
mem_k_index[4514] = 20885;
mem_k_index[4515] = 20887;
mem_k_index[4516] = 20890;
mem_k_index[4517] = 20892;
mem_k_index[4518] = 20895;
mem_k_index[4519] = 20897;
mem_k_index[4520] = 20900;
mem_k_index[4521] = 20902;
mem_k_index[4522] = 20905;
mem_k_index[4523] = 20908;
mem_k_index[4524] = 20910;
mem_k_index[4525] = 20913;
mem_k_index[4526] = 20915;
mem_k_index[4527] = 20918;
mem_k_index[4528] = 20920;
mem_k_index[4529] = 20923;
mem_k_index[4530] = 20925;
mem_k_index[4531] = 20928;
mem_k_index[4532] = 20930;
mem_k_index[4533] = 20933;
mem_k_index[4534] = 20935;
mem_k_index[4535] = 20938;
mem_k_index[4536] = 20940;
mem_k_index[4537] = 20943;
mem_k_index[4538] = 20945;
mem_k_index[4539] = 20948;
mem_k_index[4540] = 20950;
mem_k_index[4541] = 20953;
mem_k_index[4542] = 20955;
mem_k_index[4543] = 20958;
mem_k_index[4544] = 20960;
mem_k_index[4545] = 20963;
mem_k_index[4546] = 20965;
mem_k_index[4547] = 20968;
mem_k_index[4548] = 20970;
mem_k_index[4549] = 20973;
mem_k_index[4550] = 20975;
mem_k_index[4551] = 20978;
mem_k_index[4552] = 20980;
mem_k_index[4553] = 20983;
mem_k_index[4554] = 20985;
mem_k_index[4555] = 20988;
mem_k_index[4556] = 20990;
mem_k_index[4557] = 20993;
mem_k_index[4558] = 20995;
mem_k_index[4559] = 20998;
mem_k_index[4560] = 21000;
mem_k_index[4561] = 21003;
mem_k_index[4562] = 21005;
mem_k_index[4563] = 21008;
mem_k_index[4564] = 21010;
mem_k_index[4565] = 21013;
mem_k_index[4566] = 21016;
mem_k_index[4567] = 21018;
mem_k_index[4568] = 21021;
mem_k_index[4569] = 21023;
mem_k_index[4570] = 21026;
mem_k_index[4571] = 21028;
mem_k_index[4572] = 21031;
mem_k_index[4573] = 21033;
mem_k_index[4574] = 21036;
mem_k_index[4575] = 21038;
mem_k_index[4576] = 21041;
mem_k_index[4577] = 21043;
mem_k_index[4578] = 21046;
mem_k_index[4579] = 21048;
mem_k_index[4580] = 21051;
mem_k_index[4581] = 21053;
mem_k_index[4582] = 21056;
mem_k_index[4583] = 21058;
mem_k_index[4584] = 21061;
mem_k_index[4585] = 21063;
mem_k_index[4586] = 21066;
mem_k_index[4587] = 21068;
mem_k_index[4588] = 21071;
mem_k_index[4589] = 21073;
mem_k_index[4590] = 21076;
mem_k_index[4591] = 21078;
mem_k_index[4592] = 21081;
mem_k_index[4593] = 21083;
mem_k_index[4594] = 21086;
mem_k_index[4595] = 21088;
mem_k_index[4596] = 21091;
mem_k_index[4597] = 21093;
mem_k_index[4598] = 21096;
mem_k_index[4599] = 21098;
mem_k_index[4600] = 21101;
mem_k_index[4601] = 21103;
mem_k_index[4602] = 21106;
mem_k_index[4603] = 21108;
mem_k_index[4604] = 21111;
mem_k_index[4605] = 21113;
mem_k_index[4606] = 21116;
mem_k_index[4607] = 21118;
mem_k_index[4608] = 21440;
mem_k_index[4609] = 21442;
mem_k_index[4610] = 21445;
mem_k_index[4611] = 21447;
mem_k_index[4612] = 21450;
mem_k_index[4613] = 21452;
mem_k_index[4614] = 21455;
mem_k_index[4615] = 21457;
mem_k_index[4616] = 21460;
mem_k_index[4617] = 21462;
mem_k_index[4618] = 21465;
mem_k_index[4619] = 21467;
mem_k_index[4620] = 21470;
mem_k_index[4621] = 21472;
mem_k_index[4622] = 21475;
mem_k_index[4623] = 21477;
mem_k_index[4624] = 21480;
mem_k_index[4625] = 21482;
mem_k_index[4626] = 21485;
mem_k_index[4627] = 21487;
mem_k_index[4628] = 21490;
mem_k_index[4629] = 21492;
mem_k_index[4630] = 21495;
mem_k_index[4631] = 21497;
mem_k_index[4632] = 21500;
mem_k_index[4633] = 21502;
mem_k_index[4634] = 21505;
mem_k_index[4635] = 21507;
mem_k_index[4636] = 21510;
mem_k_index[4637] = 21512;
mem_k_index[4638] = 21515;
mem_k_index[4639] = 21517;
mem_k_index[4640] = 21520;
mem_k_index[4641] = 21522;
mem_k_index[4642] = 21525;
mem_k_index[4643] = 21527;
mem_k_index[4644] = 21530;
mem_k_index[4645] = 21532;
mem_k_index[4646] = 21535;
mem_k_index[4647] = 21537;
mem_k_index[4648] = 21540;
mem_k_index[4649] = 21542;
mem_k_index[4650] = 21545;
mem_k_index[4651] = 21548;
mem_k_index[4652] = 21550;
mem_k_index[4653] = 21553;
mem_k_index[4654] = 21555;
mem_k_index[4655] = 21558;
mem_k_index[4656] = 21560;
mem_k_index[4657] = 21563;
mem_k_index[4658] = 21565;
mem_k_index[4659] = 21568;
mem_k_index[4660] = 21570;
mem_k_index[4661] = 21573;
mem_k_index[4662] = 21575;
mem_k_index[4663] = 21578;
mem_k_index[4664] = 21580;
mem_k_index[4665] = 21583;
mem_k_index[4666] = 21585;
mem_k_index[4667] = 21588;
mem_k_index[4668] = 21590;
mem_k_index[4669] = 21593;
mem_k_index[4670] = 21595;
mem_k_index[4671] = 21598;
mem_k_index[4672] = 21600;
mem_k_index[4673] = 21603;
mem_k_index[4674] = 21605;
mem_k_index[4675] = 21608;
mem_k_index[4676] = 21610;
mem_k_index[4677] = 21613;
mem_k_index[4678] = 21615;
mem_k_index[4679] = 21618;
mem_k_index[4680] = 21620;
mem_k_index[4681] = 21623;
mem_k_index[4682] = 21625;
mem_k_index[4683] = 21628;
mem_k_index[4684] = 21630;
mem_k_index[4685] = 21633;
mem_k_index[4686] = 21635;
mem_k_index[4687] = 21638;
mem_k_index[4688] = 21640;
mem_k_index[4689] = 21643;
mem_k_index[4690] = 21645;
mem_k_index[4691] = 21648;
mem_k_index[4692] = 21650;
mem_k_index[4693] = 21653;
mem_k_index[4694] = 21656;
mem_k_index[4695] = 21658;
mem_k_index[4696] = 21661;
mem_k_index[4697] = 21663;
mem_k_index[4698] = 21666;
mem_k_index[4699] = 21668;
mem_k_index[4700] = 21671;
mem_k_index[4701] = 21673;
mem_k_index[4702] = 21676;
mem_k_index[4703] = 21678;
mem_k_index[4704] = 21681;
mem_k_index[4705] = 21683;
mem_k_index[4706] = 21686;
mem_k_index[4707] = 21688;
mem_k_index[4708] = 21691;
mem_k_index[4709] = 21693;
mem_k_index[4710] = 21696;
mem_k_index[4711] = 21698;
mem_k_index[4712] = 21701;
mem_k_index[4713] = 21703;
mem_k_index[4714] = 21706;
mem_k_index[4715] = 21708;
mem_k_index[4716] = 21711;
mem_k_index[4717] = 21713;
mem_k_index[4718] = 21716;
mem_k_index[4719] = 21718;
mem_k_index[4720] = 21721;
mem_k_index[4721] = 21723;
mem_k_index[4722] = 21726;
mem_k_index[4723] = 21728;
mem_k_index[4724] = 21731;
mem_k_index[4725] = 21733;
mem_k_index[4726] = 21736;
mem_k_index[4727] = 21738;
mem_k_index[4728] = 21741;
mem_k_index[4729] = 21743;
mem_k_index[4730] = 21746;
mem_k_index[4731] = 21748;
mem_k_index[4732] = 21751;
mem_k_index[4733] = 21753;
mem_k_index[4734] = 21756;
mem_k_index[4735] = 21758;
mem_k_index[4736] = 22080;
mem_k_index[4737] = 22082;
mem_k_index[4738] = 22085;
mem_k_index[4739] = 22087;
mem_k_index[4740] = 22090;
mem_k_index[4741] = 22092;
mem_k_index[4742] = 22095;
mem_k_index[4743] = 22097;
mem_k_index[4744] = 22100;
mem_k_index[4745] = 22102;
mem_k_index[4746] = 22105;
mem_k_index[4747] = 22107;
mem_k_index[4748] = 22110;
mem_k_index[4749] = 22112;
mem_k_index[4750] = 22115;
mem_k_index[4751] = 22117;
mem_k_index[4752] = 22120;
mem_k_index[4753] = 22122;
mem_k_index[4754] = 22125;
mem_k_index[4755] = 22127;
mem_k_index[4756] = 22130;
mem_k_index[4757] = 22132;
mem_k_index[4758] = 22135;
mem_k_index[4759] = 22137;
mem_k_index[4760] = 22140;
mem_k_index[4761] = 22142;
mem_k_index[4762] = 22145;
mem_k_index[4763] = 22147;
mem_k_index[4764] = 22150;
mem_k_index[4765] = 22152;
mem_k_index[4766] = 22155;
mem_k_index[4767] = 22157;
mem_k_index[4768] = 22160;
mem_k_index[4769] = 22162;
mem_k_index[4770] = 22165;
mem_k_index[4771] = 22167;
mem_k_index[4772] = 22170;
mem_k_index[4773] = 22172;
mem_k_index[4774] = 22175;
mem_k_index[4775] = 22177;
mem_k_index[4776] = 22180;
mem_k_index[4777] = 22182;
mem_k_index[4778] = 22185;
mem_k_index[4779] = 22188;
mem_k_index[4780] = 22190;
mem_k_index[4781] = 22193;
mem_k_index[4782] = 22195;
mem_k_index[4783] = 22198;
mem_k_index[4784] = 22200;
mem_k_index[4785] = 22203;
mem_k_index[4786] = 22205;
mem_k_index[4787] = 22208;
mem_k_index[4788] = 22210;
mem_k_index[4789] = 22213;
mem_k_index[4790] = 22215;
mem_k_index[4791] = 22218;
mem_k_index[4792] = 22220;
mem_k_index[4793] = 22223;
mem_k_index[4794] = 22225;
mem_k_index[4795] = 22228;
mem_k_index[4796] = 22230;
mem_k_index[4797] = 22233;
mem_k_index[4798] = 22235;
mem_k_index[4799] = 22238;
mem_k_index[4800] = 22240;
mem_k_index[4801] = 22243;
mem_k_index[4802] = 22245;
mem_k_index[4803] = 22248;
mem_k_index[4804] = 22250;
mem_k_index[4805] = 22253;
mem_k_index[4806] = 22255;
mem_k_index[4807] = 22258;
mem_k_index[4808] = 22260;
mem_k_index[4809] = 22263;
mem_k_index[4810] = 22265;
mem_k_index[4811] = 22268;
mem_k_index[4812] = 22270;
mem_k_index[4813] = 22273;
mem_k_index[4814] = 22275;
mem_k_index[4815] = 22278;
mem_k_index[4816] = 22280;
mem_k_index[4817] = 22283;
mem_k_index[4818] = 22285;
mem_k_index[4819] = 22288;
mem_k_index[4820] = 22290;
mem_k_index[4821] = 22293;
mem_k_index[4822] = 22296;
mem_k_index[4823] = 22298;
mem_k_index[4824] = 22301;
mem_k_index[4825] = 22303;
mem_k_index[4826] = 22306;
mem_k_index[4827] = 22308;
mem_k_index[4828] = 22311;
mem_k_index[4829] = 22313;
mem_k_index[4830] = 22316;
mem_k_index[4831] = 22318;
mem_k_index[4832] = 22321;
mem_k_index[4833] = 22323;
mem_k_index[4834] = 22326;
mem_k_index[4835] = 22328;
mem_k_index[4836] = 22331;
mem_k_index[4837] = 22333;
mem_k_index[4838] = 22336;
mem_k_index[4839] = 22338;
mem_k_index[4840] = 22341;
mem_k_index[4841] = 22343;
mem_k_index[4842] = 22346;
mem_k_index[4843] = 22348;
mem_k_index[4844] = 22351;
mem_k_index[4845] = 22353;
mem_k_index[4846] = 22356;
mem_k_index[4847] = 22358;
mem_k_index[4848] = 22361;
mem_k_index[4849] = 22363;
mem_k_index[4850] = 22366;
mem_k_index[4851] = 22368;
mem_k_index[4852] = 22371;
mem_k_index[4853] = 22373;
mem_k_index[4854] = 22376;
mem_k_index[4855] = 22378;
mem_k_index[4856] = 22381;
mem_k_index[4857] = 22383;
mem_k_index[4858] = 22386;
mem_k_index[4859] = 22388;
mem_k_index[4860] = 22391;
mem_k_index[4861] = 22393;
mem_k_index[4862] = 22396;
mem_k_index[4863] = 22398;
mem_k_index[4864] = 22720;
mem_k_index[4865] = 22722;
mem_k_index[4866] = 22725;
mem_k_index[4867] = 22727;
mem_k_index[4868] = 22730;
mem_k_index[4869] = 22732;
mem_k_index[4870] = 22735;
mem_k_index[4871] = 22737;
mem_k_index[4872] = 22740;
mem_k_index[4873] = 22742;
mem_k_index[4874] = 22745;
mem_k_index[4875] = 22747;
mem_k_index[4876] = 22750;
mem_k_index[4877] = 22752;
mem_k_index[4878] = 22755;
mem_k_index[4879] = 22757;
mem_k_index[4880] = 22760;
mem_k_index[4881] = 22762;
mem_k_index[4882] = 22765;
mem_k_index[4883] = 22767;
mem_k_index[4884] = 22770;
mem_k_index[4885] = 22772;
mem_k_index[4886] = 22775;
mem_k_index[4887] = 22777;
mem_k_index[4888] = 22780;
mem_k_index[4889] = 22782;
mem_k_index[4890] = 22785;
mem_k_index[4891] = 22787;
mem_k_index[4892] = 22790;
mem_k_index[4893] = 22792;
mem_k_index[4894] = 22795;
mem_k_index[4895] = 22797;
mem_k_index[4896] = 22800;
mem_k_index[4897] = 22802;
mem_k_index[4898] = 22805;
mem_k_index[4899] = 22807;
mem_k_index[4900] = 22810;
mem_k_index[4901] = 22812;
mem_k_index[4902] = 22815;
mem_k_index[4903] = 22817;
mem_k_index[4904] = 22820;
mem_k_index[4905] = 22822;
mem_k_index[4906] = 22825;
mem_k_index[4907] = 22828;
mem_k_index[4908] = 22830;
mem_k_index[4909] = 22833;
mem_k_index[4910] = 22835;
mem_k_index[4911] = 22838;
mem_k_index[4912] = 22840;
mem_k_index[4913] = 22843;
mem_k_index[4914] = 22845;
mem_k_index[4915] = 22848;
mem_k_index[4916] = 22850;
mem_k_index[4917] = 22853;
mem_k_index[4918] = 22855;
mem_k_index[4919] = 22858;
mem_k_index[4920] = 22860;
mem_k_index[4921] = 22863;
mem_k_index[4922] = 22865;
mem_k_index[4923] = 22868;
mem_k_index[4924] = 22870;
mem_k_index[4925] = 22873;
mem_k_index[4926] = 22875;
mem_k_index[4927] = 22878;
mem_k_index[4928] = 22880;
mem_k_index[4929] = 22883;
mem_k_index[4930] = 22885;
mem_k_index[4931] = 22888;
mem_k_index[4932] = 22890;
mem_k_index[4933] = 22893;
mem_k_index[4934] = 22895;
mem_k_index[4935] = 22898;
mem_k_index[4936] = 22900;
mem_k_index[4937] = 22903;
mem_k_index[4938] = 22905;
mem_k_index[4939] = 22908;
mem_k_index[4940] = 22910;
mem_k_index[4941] = 22913;
mem_k_index[4942] = 22915;
mem_k_index[4943] = 22918;
mem_k_index[4944] = 22920;
mem_k_index[4945] = 22923;
mem_k_index[4946] = 22925;
mem_k_index[4947] = 22928;
mem_k_index[4948] = 22930;
mem_k_index[4949] = 22933;
mem_k_index[4950] = 22936;
mem_k_index[4951] = 22938;
mem_k_index[4952] = 22941;
mem_k_index[4953] = 22943;
mem_k_index[4954] = 22946;
mem_k_index[4955] = 22948;
mem_k_index[4956] = 22951;
mem_k_index[4957] = 22953;
mem_k_index[4958] = 22956;
mem_k_index[4959] = 22958;
mem_k_index[4960] = 22961;
mem_k_index[4961] = 22963;
mem_k_index[4962] = 22966;
mem_k_index[4963] = 22968;
mem_k_index[4964] = 22971;
mem_k_index[4965] = 22973;
mem_k_index[4966] = 22976;
mem_k_index[4967] = 22978;
mem_k_index[4968] = 22981;
mem_k_index[4969] = 22983;
mem_k_index[4970] = 22986;
mem_k_index[4971] = 22988;
mem_k_index[4972] = 22991;
mem_k_index[4973] = 22993;
mem_k_index[4974] = 22996;
mem_k_index[4975] = 22998;
mem_k_index[4976] = 23001;
mem_k_index[4977] = 23003;
mem_k_index[4978] = 23006;
mem_k_index[4979] = 23008;
mem_k_index[4980] = 23011;
mem_k_index[4981] = 23013;
mem_k_index[4982] = 23016;
mem_k_index[4983] = 23018;
mem_k_index[4984] = 23021;
mem_k_index[4985] = 23023;
mem_k_index[4986] = 23026;
mem_k_index[4987] = 23028;
mem_k_index[4988] = 23031;
mem_k_index[4989] = 23033;
mem_k_index[4990] = 23036;
mem_k_index[4991] = 23038;
mem_k_index[4992] = 23360;
mem_k_index[4993] = 23362;
mem_k_index[4994] = 23365;
mem_k_index[4995] = 23367;
mem_k_index[4996] = 23370;
mem_k_index[4997] = 23372;
mem_k_index[4998] = 23375;
mem_k_index[4999] = 23377;
mem_k_index[5000] = 23380;
mem_k_index[5001] = 23382;
mem_k_index[5002] = 23385;
mem_k_index[5003] = 23387;
mem_k_index[5004] = 23390;
mem_k_index[5005] = 23392;
mem_k_index[5006] = 23395;
mem_k_index[5007] = 23397;
mem_k_index[5008] = 23400;
mem_k_index[5009] = 23402;
mem_k_index[5010] = 23405;
mem_k_index[5011] = 23407;
mem_k_index[5012] = 23410;
mem_k_index[5013] = 23412;
mem_k_index[5014] = 23415;
mem_k_index[5015] = 23417;
mem_k_index[5016] = 23420;
mem_k_index[5017] = 23422;
mem_k_index[5018] = 23425;
mem_k_index[5019] = 23427;
mem_k_index[5020] = 23430;
mem_k_index[5021] = 23432;
mem_k_index[5022] = 23435;
mem_k_index[5023] = 23437;
mem_k_index[5024] = 23440;
mem_k_index[5025] = 23442;
mem_k_index[5026] = 23445;
mem_k_index[5027] = 23447;
mem_k_index[5028] = 23450;
mem_k_index[5029] = 23452;
mem_k_index[5030] = 23455;
mem_k_index[5031] = 23457;
mem_k_index[5032] = 23460;
mem_k_index[5033] = 23462;
mem_k_index[5034] = 23465;
mem_k_index[5035] = 23468;
mem_k_index[5036] = 23470;
mem_k_index[5037] = 23473;
mem_k_index[5038] = 23475;
mem_k_index[5039] = 23478;
mem_k_index[5040] = 23480;
mem_k_index[5041] = 23483;
mem_k_index[5042] = 23485;
mem_k_index[5043] = 23488;
mem_k_index[5044] = 23490;
mem_k_index[5045] = 23493;
mem_k_index[5046] = 23495;
mem_k_index[5047] = 23498;
mem_k_index[5048] = 23500;
mem_k_index[5049] = 23503;
mem_k_index[5050] = 23505;
mem_k_index[5051] = 23508;
mem_k_index[5052] = 23510;
mem_k_index[5053] = 23513;
mem_k_index[5054] = 23515;
mem_k_index[5055] = 23518;
mem_k_index[5056] = 23520;
mem_k_index[5057] = 23523;
mem_k_index[5058] = 23525;
mem_k_index[5059] = 23528;
mem_k_index[5060] = 23530;
mem_k_index[5061] = 23533;
mem_k_index[5062] = 23535;
mem_k_index[5063] = 23538;
mem_k_index[5064] = 23540;
mem_k_index[5065] = 23543;
mem_k_index[5066] = 23545;
mem_k_index[5067] = 23548;
mem_k_index[5068] = 23550;
mem_k_index[5069] = 23553;
mem_k_index[5070] = 23555;
mem_k_index[5071] = 23558;
mem_k_index[5072] = 23560;
mem_k_index[5073] = 23563;
mem_k_index[5074] = 23565;
mem_k_index[5075] = 23568;
mem_k_index[5076] = 23570;
mem_k_index[5077] = 23573;
mem_k_index[5078] = 23576;
mem_k_index[5079] = 23578;
mem_k_index[5080] = 23581;
mem_k_index[5081] = 23583;
mem_k_index[5082] = 23586;
mem_k_index[5083] = 23588;
mem_k_index[5084] = 23591;
mem_k_index[5085] = 23593;
mem_k_index[5086] = 23596;
mem_k_index[5087] = 23598;
mem_k_index[5088] = 23601;
mem_k_index[5089] = 23603;
mem_k_index[5090] = 23606;
mem_k_index[5091] = 23608;
mem_k_index[5092] = 23611;
mem_k_index[5093] = 23613;
mem_k_index[5094] = 23616;
mem_k_index[5095] = 23618;
mem_k_index[5096] = 23621;
mem_k_index[5097] = 23623;
mem_k_index[5098] = 23626;
mem_k_index[5099] = 23628;
mem_k_index[5100] = 23631;
mem_k_index[5101] = 23633;
mem_k_index[5102] = 23636;
mem_k_index[5103] = 23638;
mem_k_index[5104] = 23641;
mem_k_index[5105] = 23643;
mem_k_index[5106] = 23646;
mem_k_index[5107] = 23648;
mem_k_index[5108] = 23651;
mem_k_index[5109] = 23653;
mem_k_index[5110] = 23656;
mem_k_index[5111] = 23658;
mem_k_index[5112] = 23661;
mem_k_index[5113] = 23663;
mem_k_index[5114] = 23666;
mem_k_index[5115] = 23668;
mem_k_index[5116] = 23671;
mem_k_index[5117] = 23673;
mem_k_index[5118] = 23676;
mem_k_index[5119] = 23678;
mem_k_index[5120] = 24000;
mem_k_index[5121] = 24002;
mem_k_index[5122] = 24005;
mem_k_index[5123] = 24007;
mem_k_index[5124] = 24010;
mem_k_index[5125] = 24012;
mem_k_index[5126] = 24015;
mem_k_index[5127] = 24017;
mem_k_index[5128] = 24020;
mem_k_index[5129] = 24022;
mem_k_index[5130] = 24025;
mem_k_index[5131] = 24027;
mem_k_index[5132] = 24030;
mem_k_index[5133] = 24032;
mem_k_index[5134] = 24035;
mem_k_index[5135] = 24037;
mem_k_index[5136] = 24040;
mem_k_index[5137] = 24042;
mem_k_index[5138] = 24045;
mem_k_index[5139] = 24047;
mem_k_index[5140] = 24050;
mem_k_index[5141] = 24052;
mem_k_index[5142] = 24055;
mem_k_index[5143] = 24057;
mem_k_index[5144] = 24060;
mem_k_index[5145] = 24062;
mem_k_index[5146] = 24065;
mem_k_index[5147] = 24067;
mem_k_index[5148] = 24070;
mem_k_index[5149] = 24072;
mem_k_index[5150] = 24075;
mem_k_index[5151] = 24077;
mem_k_index[5152] = 24080;
mem_k_index[5153] = 24082;
mem_k_index[5154] = 24085;
mem_k_index[5155] = 24087;
mem_k_index[5156] = 24090;
mem_k_index[5157] = 24092;
mem_k_index[5158] = 24095;
mem_k_index[5159] = 24097;
mem_k_index[5160] = 24100;
mem_k_index[5161] = 24102;
mem_k_index[5162] = 24105;
mem_k_index[5163] = 24108;
mem_k_index[5164] = 24110;
mem_k_index[5165] = 24113;
mem_k_index[5166] = 24115;
mem_k_index[5167] = 24118;
mem_k_index[5168] = 24120;
mem_k_index[5169] = 24123;
mem_k_index[5170] = 24125;
mem_k_index[5171] = 24128;
mem_k_index[5172] = 24130;
mem_k_index[5173] = 24133;
mem_k_index[5174] = 24135;
mem_k_index[5175] = 24138;
mem_k_index[5176] = 24140;
mem_k_index[5177] = 24143;
mem_k_index[5178] = 24145;
mem_k_index[5179] = 24148;
mem_k_index[5180] = 24150;
mem_k_index[5181] = 24153;
mem_k_index[5182] = 24155;
mem_k_index[5183] = 24158;
mem_k_index[5184] = 24160;
mem_k_index[5185] = 24163;
mem_k_index[5186] = 24165;
mem_k_index[5187] = 24168;
mem_k_index[5188] = 24170;
mem_k_index[5189] = 24173;
mem_k_index[5190] = 24175;
mem_k_index[5191] = 24178;
mem_k_index[5192] = 24180;
mem_k_index[5193] = 24183;
mem_k_index[5194] = 24185;
mem_k_index[5195] = 24188;
mem_k_index[5196] = 24190;
mem_k_index[5197] = 24193;
mem_k_index[5198] = 24195;
mem_k_index[5199] = 24198;
mem_k_index[5200] = 24200;
mem_k_index[5201] = 24203;
mem_k_index[5202] = 24205;
mem_k_index[5203] = 24208;
mem_k_index[5204] = 24210;
mem_k_index[5205] = 24213;
mem_k_index[5206] = 24216;
mem_k_index[5207] = 24218;
mem_k_index[5208] = 24221;
mem_k_index[5209] = 24223;
mem_k_index[5210] = 24226;
mem_k_index[5211] = 24228;
mem_k_index[5212] = 24231;
mem_k_index[5213] = 24233;
mem_k_index[5214] = 24236;
mem_k_index[5215] = 24238;
mem_k_index[5216] = 24241;
mem_k_index[5217] = 24243;
mem_k_index[5218] = 24246;
mem_k_index[5219] = 24248;
mem_k_index[5220] = 24251;
mem_k_index[5221] = 24253;
mem_k_index[5222] = 24256;
mem_k_index[5223] = 24258;
mem_k_index[5224] = 24261;
mem_k_index[5225] = 24263;
mem_k_index[5226] = 24266;
mem_k_index[5227] = 24268;
mem_k_index[5228] = 24271;
mem_k_index[5229] = 24273;
mem_k_index[5230] = 24276;
mem_k_index[5231] = 24278;
mem_k_index[5232] = 24281;
mem_k_index[5233] = 24283;
mem_k_index[5234] = 24286;
mem_k_index[5235] = 24288;
mem_k_index[5236] = 24291;
mem_k_index[5237] = 24293;
mem_k_index[5238] = 24296;
mem_k_index[5239] = 24298;
mem_k_index[5240] = 24301;
mem_k_index[5241] = 24303;
mem_k_index[5242] = 24306;
mem_k_index[5243] = 24308;
mem_k_index[5244] = 24311;
mem_k_index[5245] = 24313;
mem_k_index[5246] = 24316;
mem_k_index[5247] = 24318;
mem_k_index[5248] = 24640;
mem_k_index[5249] = 24642;
mem_k_index[5250] = 24645;
mem_k_index[5251] = 24647;
mem_k_index[5252] = 24650;
mem_k_index[5253] = 24652;
mem_k_index[5254] = 24655;
mem_k_index[5255] = 24657;
mem_k_index[5256] = 24660;
mem_k_index[5257] = 24662;
mem_k_index[5258] = 24665;
mem_k_index[5259] = 24667;
mem_k_index[5260] = 24670;
mem_k_index[5261] = 24672;
mem_k_index[5262] = 24675;
mem_k_index[5263] = 24677;
mem_k_index[5264] = 24680;
mem_k_index[5265] = 24682;
mem_k_index[5266] = 24685;
mem_k_index[5267] = 24687;
mem_k_index[5268] = 24690;
mem_k_index[5269] = 24692;
mem_k_index[5270] = 24695;
mem_k_index[5271] = 24697;
mem_k_index[5272] = 24700;
mem_k_index[5273] = 24702;
mem_k_index[5274] = 24705;
mem_k_index[5275] = 24707;
mem_k_index[5276] = 24710;
mem_k_index[5277] = 24712;
mem_k_index[5278] = 24715;
mem_k_index[5279] = 24717;
mem_k_index[5280] = 24720;
mem_k_index[5281] = 24722;
mem_k_index[5282] = 24725;
mem_k_index[5283] = 24727;
mem_k_index[5284] = 24730;
mem_k_index[5285] = 24732;
mem_k_index[5286] = 24735;
mem_k_index[5287] = 24737;
mem_k_index[5288] = 24740;
mem_k_index[5289] = 24742;
mem_k_index[5290] = 24745;
mem_k_index[5291] = 24748;
mem_k_index[5292] = 24750;
mem_k_index[5293] = 24753;
mem_k_index[5294] = 24755;
mem_k_index[5295] = 24758;
mem_k_index[5296] = 24760;
mem_k_index[5297] = 24763;
mem_k_index[5298] = 24765;
mem_k_index[5299] = 24768;
mem_k_index[5300] = 24770;
mem_k_index[5301] = 24773;
mem_k_index[5302] = 24775;
mem_k_index[5303] = 24778;
mem_k_index[5304] = 24780;
mem_k_index[5305] = 24783;
mem_k_index[5306] = 24785;
mem_k_index[5307] = 24788;
mem_k_index[5308] = 24790;
mem_k_index[5309] = 24793;
mem_k_index[5310] = 24795;
mem_k_index[5311] = 24798;
mem_k_index[5312] = 24800;
mem_k_index[5313] = 24803;
mem_k_index[5314] = 24805;
mem_k_index[5315] = 24808;
mem_k_index[5316] = 24810;
mem_k_index[5317] = 24813;
mem_k_index[5318] = 24815;
mem_k_index[5319] = 24818;
mem_k_index[5320] = 24820;
mem_k_index[5321] = 24823;
mem_k_index[5322] = 24825;
mem_k_index[5323] = 24828;
mem_k_index[5324] = 24830;
mem_k_index[5325] = 24833;
mem_k_index[5326] = 24835;
mem_k_index[5327] = 24838;
mem_k_index[5328] = 24840;
mem_k_index[5329] = 24843;
mem_k_index[5330] = 24845;
mem_k_index[5331] = 24848;
mem_k_index[5332] = 24850;
mem_k_index[5333] = 24853;
mem_k_index[5334] = 24856;
mem_k_index[5335] = 24858;
mem_k_index[5336] = 24861;
mem_k_index[5337] = 24863;
mem_k_index[5338] = 24866;
mem_k_index[5339] = 24868;
mem_k_index[5340] = 24871;
mem_k_index[5341] = 24873;
mem_k_index[5342] = 24876;
mem_k_index[5343] = 24878;
mem_k_index[5344] = 24881;
mem_k_index[5345] = 24883;
mem_k_index[5346] = 24886;
mem_k_index[5347] = 24888;
mem_k_index[5348] = 24891;
mem_k_index[5349] = 24893;
mem_k_index[5350] = 24896;
mem_k_index[5351] = 24898;
mem_k_index[5352] = 24901;
mem_k_index[5353] = 24903;
mem_k_index[5354] = 24906;
mem_k_index[5355] = 24908;
mem_k_index[5356] = 24911;
mem_k_index[5357] = 24913;
mem_k_index[5358] = 24916;
mem_k_index[5359] = 24918;
mem_k_index[5360] = 24921;
mem_k_index[5361] = 24923;
mem_k_index[5362] = 24926;
mem_k_index[5363] = 24928;
mem_k_index[5364] = 24931;
mem_k_index[5365] = 24933;
mem_k_index[5366] = 24936;
mem_k_index[5367] = 24938;
mem_k_index[5368] = 24941;
mem_k_index[5369] = 24943;
mem_k_index[5370] = 24946;
mem_k_index[5371] = 24948;
mem_k_index[5372] = 24951;
mem_k_index[5373] = 24953;
mem_k_index[5374] = 24956;
mem_k_index[5375] = 24958;
mem_k_index[5376] = 25280;
mem_k_index[5377] = 25282;
mem_k_index[5378] = 25285;
mem_k_index[5379] = 25287;
mem_k_index[5380] = 25290;
mem_k_index[5381] = 25292;
mem_k_index[5382] = 25295;
mem_k_index[5383] = 25297;
mem_k_index[5384] = 25300;
mem_k_index[5385] = 25302;
mem_k_index[5386] = 25305;
mem_k_index[5387] = 25307;
mem_k_index[5388] = 25310;
mem_k_index[5389] = 25312;
mem_k_index[5390] = 25315;
mem_k_index[5391] = 25317;
mem_k_index[5392] = 25320;
mem_k_index[5393] = 25322;
mem_k_index[5394] = 25325;
mem_k_index[5395] = 25327;
mem_k_index[5396] = 25330;
mem_k_index[5397] = 25332;
mem_k_index[5398] = 25335;
mem_k_index[5399] = 25337;
mem_k_index[5400] = 25340;
mem_k_index[5401] = 25342;
mem_k_index[5402] = 25345;
mem_k_index[5403] = 25347;
mem_k_index[5404] = 25350;
mem_k_index[5405] = 25352;
mem_k_index[5406] = 25355;
mem_k_index[5407] = 25357;
mem_k_index[5408] = 25360;
mem_k_index[5409] = 25362;
mem_k_index[5410] = 25365;
mem_k_index[5411] = 25367;
mem_k_index[5412] = 25370;
mem_k_index[5413] = 25372;
mem_k_index[5414] = 25375;
mem_k_index[5415] = 25377;
mem_k_index[5416] = 25380;
mem_k_index[5417] = 25382;
mem_k_index[5418] = 25385;
mem_k_index[5419] = 25388;
mem_k_index[5420] = 25390;
mem_k_index[5421] = 25393;
mem_k_index[5422] = 25395;
mem_k_index[5423] = 25398;
mem_k_index[5424] = 25400;
mem_k_index[5425] = 25403;
mem_k_index[5426] = 25405;
mem_k_index[5427] = 25408;
mem_k_index[5428] = 25410;
mem_k_index[5429] = 25413;
mem_k_index[5430] = 25415;
mem_k_index[5431] = 25418;
mem_k_index[5432] = 25420;
mem_k_index[5433] = 25423;
mem_k_index[5434] = 25425;
mem_k_index[5435] = 25428;
mem_k_index[5436] = 25430;
mem_k_index[5437] = 25433;
mem_k_index[5438] = 25435;
mem_k_index[5439] = 25438;
mem_k_index[5440] = 25440;
mem_k_index[5441] = 25443;
mem_k_index[5442] = 25445;
mem_k_index[5443] = 25448;
mem_k_index[5444] = 25450;
mem_k_index[5445] = 25453;
mem_k_index[5446] = 25455;
mem_k_index[5447] = 25458;
mem_k_index[5448] = 25460;
mem_k_index[5449] = 25463;
mem_k_index[5450] = 25465;
mem_k_index[5451] = 25468;
mem_k_index[5452] = 25470;
mem_k_index[5453] = 25473;
mem_k_index[5454] = 25475;
mem_k_index[5455] = 25478;
mem_k_index[5456] = 25480;
mem_k_index[5457] = 25483;
mem_k_index[5458] = 25485;
mem_k_index[5459] = 25488;
mem_k_index[5460] = 25490;
mem_k_index[5461] = 25493;
mem_k_index[5462] = 25496;
mem_k_index[5463] = 25498;
mem_k_index[5464] = 25501;
mem_k_index[5465] = 25503;
mem_k_index[5466] = 25506;
mem_k_index[5467] = 25508;
mem_k_index[5468] = 25511;
mem_k_index[5469] = 25513;
mem_k_index[5470] = 25516;
mem_k_index[5471] = 25518;
mem_k_index[5472] = 25521;
mem_k_index[5473] = 25523;
mem_k_index[5474] = 25526;
mem_k_index[5475] = 25528;
mem_k_index[5476] = 25531;
mem_k_index[5477] = 25533;
mem_k_index[5478] = 25536;
mem_k_index[5479] = 25538;
mem_k_index[5480] = 25541;
mem_k_index[5481] = 25543;
mem_k_index[5482] = 25546;
mem_k_index[5483] = 25548;
mem_k_index[5484] = 25551;
mem_k_index[5485] = 25553;
mem_k_index[5486] = 25556;
mem_k_index[5487] = 25558;
mem_k_index[5488] = 25561;
mem_k_index[5489] = 25563;
mem_k_index[5490] = 25566;
mem_k_index[5491] = 25568;
mem_k_index[5492] = 25571;
mem_k_index[5493] = 25573;
mem_k_index[5494] = 25576;
mem_k_index[5495] = 25578;
mem_k_index[5496] = 25581;
mem_k_index[5497] = 25583;
mem_k_index[5498] = 25586;
mem_k_index[5499] = 25588;
mem_k_index[5500] = 25591;
mem_k_index[5501] = 25593;
mem_k_index[5502] = 25596;
mem_k_index[5503] = 25598;
mem_k_index[5504] = 25600;
mem_k_index[5505] = 25602;
mem_k_index[5506] = 25605;
mem_k_index[5507] = 25607;
mem_k_index[5508] = 25610;
mem_k_index[5509] = 25612;
mem_k_index[5510] = 25615;
mem_k_index[5511] = 25617;
mem_k_index[5512] = 25620;
mem_k_index[5513] = 25622;
mem_k_index[5514] = 25625;
mem_k_index[5515] = 25627;
mem_k_index[5516] = 25630;
mem_k_index[5517] = 25632;
mem_k_index[5518] = 25635;
mem_k_index[5519] = 25637;
mem_k_index[5520] = 25640;
mem_k_index[5521] = 25642;
mem_k_index[5522] = 25645;
mem_k_index[5523] = 25647;
mem_k_index[5524] = 25650;
mem_k_index[5525] = 25652;
mem_k_index[5526] = 25655;
mem_k_index[5527] = 25657;
mem_k_index[5528] = 25660;
mem_k_index[5529] = 25662;
mem_k_index[5530] = 25665;
mem_k_index[5531] = 25667;
mem_k_index[5532] = 25670;
mem_k_index[5533] = 25672;
mem_k_index[5534] = 25675;
mem_k_index[5535] = 25677;
mem_k_index[5536] = 25680;
mem_k_index[5537] = 25682;
mem_k_index[5538] = 25685;
mem_k_index[5539] = 25687;
mem_k_index[5540] = 25690;
mem_k_index[5541] = 25692;
mem_k_index[5542] = 25695;
mem_k_index[5543] = 25697;
mem_k_index[5544] = 25700;
mem_k_index[5545] = 25702;
mem_k_index[5546] = 25705;
mem_k_index[5547] = 25708;
mem_k_index[5548] = 25710;
mem_k_index[5549] = 25713;
mem_k_index[5550] = 25715;
mem_k_index[5551] = 25718;
mem_k_index[5552] = 25720;
mem_k_index[5553] = 25723;
mem_k_index[5554] = 25725;
mem_k_index[5555] = 25728;
mem_k_index[5556] = 25730;
mem_k_index[5557] = 25733;
mem_k_index[5558] = 25735;
mem_k_index[5559] = 25738;
mem_k_index[5560] = 25740;
mem_k_index[5561] = 25743;
mem_k_index[5562] = 25745;
mem_k_index[5563] = 25748;
mem_k_index[5564] = 25750;
mem_k_index[5565] = 25753;
mem_k_index[5566] = 25755;
mem_k_index[5567] = 25758;
mem_k_index[5568] = 25760;
mem_k_index[5569] = 25763;
mem_k_index[5570] = 25765;
mem_k_index[5571] = 25768;
mem_k_index[5572] = 25770;
mem_k_index[5573] = 25773;
mem_k_index[5574] = 25775;
mem_k_index[5575] = 25778;
mem_k_index[5576] = 25780;
mem_k_index[5577] = 25783;
mem_k_index[5578] = 25785;
mem_k_index[5579] = 25788;
mem_k_index[5580] = 25790;
mem_k_index[5581] = 25793;
mem_k_index[5582] = 25795;
mem_k_index[5583] = 25798;
mem_k_index[5584] = 25800;
mem_k_index[5585] = 25803;
mem_k_index[5586] = 25805;
mem_k_index[5587] = 25808;
mem_k_index[5588] = 25810;
mem_k_index[5589] = 25813;
mem_k_index[5590] = 25816;
mem_k_index[5591] = 25818;
mem_k_index[5592] = 25821;
mem_k_index[5593] = 25823;
mem_k_index[5594] = 25826;
mem_k_index[5595] = 25828;
mem_k_index[5596] = 25831;
mem_k_index[5597] = 25833;
mem_k_index[5598] = 25836;
mem_k_index[5599] = 25838;
mem_k_index[5600] = 25841;
mem_k_index[5601] = 25843;
mem_k_index[5602] = 25846;
mem_k_index[5603] = 25848;
mem_k_index[5604] = 25851;
mem_k_index[5605] = 25853;
mem_k_index[5606] = 25856;
mem_k_index[5607] = 25858;
mem_k_index[5608] = 25861;
mem_k_index[5609] = 25863;
mem_k_index[5610] = 25866;
mem_k_index[5611] = 25868;
mem_k_index[5612] = 25871;
mem_k_index[5613] = 25873;
mem_k_index[5614] = 25876;
mem_k_index[5615] = 25878;
mem_k_index[5616] = 25881;
mem_k_index[5617] = 25883;
mem_k_index[5618] = 25886;
mem_k_index[5619] = 25888;
mem_k_index[5620] = 25891;
mem_k_index[5621] = 25893;
mem_k_index[5622] = 25896;
mem_k_index[5623] = 25898;
mem_k_index[5624] = 25901;
mem_k_index[5625] = 25903;
mem_k_index[5626] = 25906;
mem_k_index[5627] = 25908;
mem_k_index[5628] = 25911;
mem_k_index[5629] = 25913;
mem_k_index[5630] = 25916;
mem_k_index[5631] = 25918;
mem_k_index[5632] = 26240;
mem_k_index[5633] = 26242;
mem_k_index[5634] = 26245;
mem_k_index[5635] = 26247;
mem_k_index[5636] = 26250;
mem_k_index[5637] = 26252;
mem_k_index[5638] = 26255;
mem_k_index[5639] = 26257;
mem_k_index[5640] = 26260;
mem_k_index[5641] = 26262;
mem_k_index[5642] = 26265;
mem_k_index[5643] = 26267;
mem_k_index[5644] = 26270;
mem_k_index[5645] = 26272;
mem_k_index[5646] = 26275;
mem_k_index[5647] = 26277;
mem_k_index[5648] = 26280;
mem_k_index[5649] = 26282;
mem_k_index[5650] = 26285;
mem_k_index[5651] = 26287;
mem_k_index[5652] = 26290;
mem_k_index[5653] = 26292;
mem_k_index[5654] = 26295;
mem_k_index[5655] = 26297;
mem_k_index[5656] = 26300;
mem_k_index[5657] = 26302;
mem_k_index[5658] = 26305;
mem_k_index[5659] = 26307;
mem_k_index[5660] = 26310;
mem_k_index[5661] = 26312;
mem_k_index[5662] = 26315;
mem_k_index[5663] = 26317;
mem_k_index[5664] = 26320;
mem_k_index[5665] = 26322;
mem_k_index[5666] = 26325;
mem_k_index[5667] = 26327;
mem_k_index[5668] = 26330;
mem_k_index[5669] = 26332;
mem_k_index[5670] = 26335;
mem_k_index[5671] = 26337;
mem_k_index[5672] = 26340;
mem_k_index[5673] = 26342;
mem_k_index[5674] = 26345;
mem_k_index[5675] = 26348;
mem_k_index[5676] = 26350;
mem_k_index[5677] = 26353;
mem_k_index[5678] = 26355;
mem_k_index[5679] = 26358;
mem_k_index[5680] = 26360;
mem_k_index[5681] = 26363;
mem_k_index[5682] = 26365;
mem_k_index[5683] = 26368;
mem_k_index[5684] = 26370;
mem_k_index[5685] = 26373;
mem_k_index[5686] = 26375;
mem_k_index[5687] = 26378;
mem_k_index[5688] = 26380;
mem_k_index[5689] = 26383;
mem_k_index[5690] = 26385;
mem_k_index[5691] = 26388;
mem_k_index[5692] = 26390;
mem_k_index[5693] = 26393;
mem_k_index[5694] = 26395;
mem_k_index[5695] = 26398;
mem_k_index[5696] = 26400;
mem_k_index[5697] = 26403;
mem_k_index[5698] = 26405;
mem_k_index[5699] = 26408;
mem_k_index[5700] = 26410;
mem_k_index[5701] = 26413;
mem_k_index[5702] = 26415;
mem_k_index[5703] = 26418;
mem_k_index[5704] = 26420;
mem_k_index[5705] = 26423;
mem_k_index[5706] = 26425;
mem_k_index[5707] = 26428;
mem_k_index[5708] = 26430;
mem_k_index[5709] = 26433;
mem_k_index[5710] = 26435;
mem_k_index[5711] = 26438;
mem_k_index[5712] = 26440;
mem_k_index[5713] = 26443;
mem_k_index[5714] = 26445;
mem_k_index[5715] = 26448;
mem_k_index[5716] = 26450;
mem_k_index[5717] = 26453;
mem_k_index[5718] = 26456;
mem_k_index[5719] = 26458;
mem_k_index[5720] = 26461;
mem_k_index[5721] = 26463;
mem_k_index[5722] = 26466;
mem_k_index[5723] = 26468;
mem_k_index[5724] = 26471;
mem_k_index[5725] = 26473;
mem_k_index[5726] = 26476;
mem_k_index[5727] = 26478;
mem_k_index[5728] = 26481;
mem_k_index[5729] = 26483;
mem_k_index[5730] = 26486;
mem_k_index[5731] = 26488;
mem_k_index[5732] = 26491;
mem_k_index[5733] = 26493;
mem_k_index[5734] = 26496;
mem_k_index[5735] = 26498;
mem_k_index[5736] = 26501;
mem_k_index[5737] = 26503;
mem_k_index[5738] = 26506;
mem_k_index[5739] = 26508;
mem_k_index[5740] = 26511;
mem_k_index[5741] = 26513;
mem_k_index[5742] = 26516;
mem_k_index[5743] = 26518;
mem_k_index[5744] = 26521;
mem_k_index[5745] = 26523;
mem_k_index[5746] = 26526;
mem_k_index[5747] = 26528;
mem_k_index[5748] = 26531;
mem_k_index[5749] = 26533;
mem_k_index[5750] = 26536;
mem_k_index[5751] = 26538;
mem_k_index[5752] = 26541;
mem_k_index[5753] = 26543;
mem_k_index[5754] = 26546;
mem_k_index[5755] = 26548;
mem_k_index[5756] = 26551;
mem_k_index[5757] = 26553;
mem_k_index[5758] = 26556;
mem_k_index[5759] = 26558;
mem_k_index[5760] = 26880;
mem_k_index[5761] = 26882;
mem_k_index[5762] = 26885;
mem_k_index[5763] = 26887;
mem_k_index[5764] = 26890;
mem_k_index[5765] = 26892;
mem_k_index[5766] = 26895;
mem_k_index[5767] = 26897;
mem_k_index[5768] = 26900;
mem_k_index[5769] = 26902;
mem_k_index[5770] = 26905;
mem_k_index[5771] = 26907;
mem_k_index[5772] = 26910;
mem_k_index[5773] = 26912;
mem_k_index[5774] = 26915;
mem_k_index[5775] = 26917;
mem_k_index[5776] = 26920;
mem_k_index[5777] = 26922;
mem_k_index[5778] = 26925;
mem_k_index[5779] = 26927;
mem_k_index[5780] = 26930;
mem_k_index[5781] = 26932;
mem_k_index[5782] = 26935;
mem_k_index[5783] = 26937;
mem_k_index[5784] = 26940;
mem_k_index[5785] = 26942;
mem_k_index[5786] = 26945;
mem_k_index[5787] = 26947;
mem_k_index[5788] = 26950;
mem_k_index[5789] = 26952;
mem_k_index[5790] = 26955;
mem_k_index[5791] = 26957;
mem_k_index[5792] = 26960;
mem_k_index[5793] = 26962;
mem_k_index[5794] = 26965;
mem_k_index[5795] = 26967;
mem_k_index[5796] = 26970;
mem_k_index[5797] = 26972;
mem_k_index[5798] = 26975;
mem_k_index[5799] = 26977;
mem_k_index[5800] = 26980;
mem_k_index[5801] = 26982;
mem_k_index[5802] = 26985;
mem_k_index[5803] = 26988;
mem_k_index[5804] = 26990;
mem_k_index[5805] = 26993;
mem_k_index[5806] = 26995;
mem_k_index[5807] = 26998;
mem_k_index[5808] = 27000;
mem_k_index[5809] = 27003;
mem_k_index[5810] = 27005;
mem_k_index[5811] = 27008;
mem_k_index[5812] = 27010;
mem_k_index[5813] = 27013;
mem_k_index[5814] = 27015;
mem_k_index[5815] = 27018;
mem_k_index[5816] = 27020;
mem_k_index[5817] = 27023;
mem_k_index[5818] = 27025;
mem_k_index[5819] = 27028;
mem_k_index[5820] = 27030;
mem_k_index[5821] = 27033;
mem_k_index[5822] = 27035;
mem_k_index[5823] = 27038;
mem_k_index[5824] = 27040;
mem_k_index[5825] = 27043;
mem_k_index[5826] = 27045;
mem_k_index[5827] = 27048;
mem_k_index[5828] = 27050;
mem_k_index[5829] = 27053;
mem_k_index[5830] = 27055;
mem_k_index[5831] = 27058;
mem_k_index[5832] = 27060;
mem_k_index[5833] = 27063;
mem_k_index[5834] = 27065;
mem_k_index[5835] = 27068;
mem_k_index[5836] = 27070;
mem_k_index[5837] = 27073;
mem_k_index[5838] = 27075;
mem_k_index[5839] = 27078;
mem_k_index[5840] = 27080;
mem_k_index[5841] = 27083;
mem_k_index[5842] = 27085;
mem_k_index[5843] = 27088;
mem_k_index[5844] = 27090;
mem_k_index[5845] = 27093;
mem_k_index[5846] = 27096;
mem_k_index[5847] = 27098;
mem_k_index[5848] = 27101;
mem_k_index[5849] = 27103;
mem_k_index[5850] = 27106;
mem_k_index[5851] = 27108;
mem_k_index[5852] = 27111;
mem_k_index[5853] = 27113;
mem_k_index[5854] = 27116;
mem_k_index[5855] = 27118;
mem_k_index[5856] = 27121;
mem_k_index[5857] = 27123;
mem_k_index[5858] = 27126;
mem_k_index[5859] = 27128;
mem_k_index[5860] = 27131;
mem_k_index[5861] = 27133;
mem_k_index[5862] = 27136;
mem_k_index[5863] = 27138;
mem_k_index[5864] = 27141;
mem_k_index[5865] = 27143;
mem_k_index[5866] = 27146;
mem_k_index[5867] = 27148;
mem_k_index[5868] = 27151;
mem_k_index[5869] = 27153;
mem_k_index[5870] = 27156;
mem_k_index[5871] = 27158;
mem_k_index[5872] = 27161;
mem_k_index[5873] = 27163;
mem_k_index[5874] = 27166;
mem_k_index[5875] = 27168;
mem_k_index[5876] = 27171;
mem_k_index[5877] = 27173;
mem_k_index[5878] = 27176;
mem_k_index[5879] = 27178;
mem_k_index[5880] = 27181;
mem_k_index[5881] = 27183;
mem_k_index[5882] = 27186;
mem_k_index[5883] = 27188;
mem_k_index[5884] = 27191;
mem_k_index[5885] = 27193;
mem_k_index[5886] = 27196;
mem_k_index[5887] = 27198;
mem_k_index[5888] = 27520;
mem_k_index[5889] = 27522;
mem_k_index[5890] = 27525;
mem_k_index[5891] = 27527;
mem_k_index[5892] = 27530;
mem_k_index[5893] = 27532;
mem_k_index[5894] = 27535;
mem_k_index[5895] = 27537;
mem_k_index[5896] = 27540;
mem_k_index[5897] = 27542;
mem_k_index[5898] = 27545;
mem_k_index[5899] = 27547;
mem_k_index[5900] = 27550;
mem_k_index[5901] = 27552;
mem_k_index[5902] = 27555;
mem_k_index[5903] = 27557;
mem_k_index[5904] = 27560;
mem_k_index[5905] = 27562;
mem_k_index[5906] = 27565;
mem_k_index[5907] = 27567;
mem_k_index[5908] = 27570;
mem_k_index[5909] = 27572;
mem_k_index[5910] = 27575;
mem_k_index[5911] = 27577;
mem_k_index[5912] = 27580;
mem_k_index[5913] = 27582;
mem_k_index[5914] = 27585;
mem_k_index[5915] = 27587;
mem_k_index[5916] = 27590;
mem_k_index[5917] = 27592;
mem_k_index[5918] = 27595;
mem_k_index[5919] = 27597;
mem_k_index[5920] = 27600;
mem_k_index[5921] = 27602;
mem_k_index[5922] = 27605;
mem_k_index[5923] = 27607;
mem_k_index[5924] = 27610;
mem_k_index[5925] = 27612;
mem_k_index[5926] = 27615;
mem_k_index[5927] = 27617;
mem_k_index[5928] = 27620;
mem_k_index[5929] = 27622;
mem_k_index[5930] = 27625;
mem_k_index[5931] = 27628;
mem_k_index[5932] = 27630;
mem_k_index[5933] = 27633;
mem_k_index[5934] = 27635;
mem_k_index[5935] = 27638;
mem_k_index[5936] = 27640;
mem_k_index[5937] = 27643;
mem_k_index[5938] = 27645;
mem_k_index[5939] = 27648;
mem_k_index[5940] = 27650;
mem_k_index[5941] = 27653;
mem_k_index[5942] = 27655;
mem_k_index[5943] = 27658;
mem_k_index[5944] = 27660;
mem_k_index[5945] = 27663;
mem_k_index[5946] = 27665;
mem_k_index[5947] = 27668;
mem_k_index[5948] = 27670;
mem_k_index[5949] = 27673;
mem_k_index[5950] = 27675;
mem_k_index[5951] = 27678;
mem_k_index[5952] = 27680;
mem_k_index[5953] = 27683;
mem_k_index[5954] = 27685;
mem_k_index[5955] = 27688;
mem_k_index[5956] = 27690;
mem_k_index[5957] = 27693;
mem_k_index[5958] = 27695;
mem_k_index[5959] = 27698;
mem_k_index[5960] = 27700;
mem_k_index[5961] = 27703;
mem_k_index[5962] = 27705;
mem_k_index[5963] = 27708;
mem_k_index[5964] = 27710;
mem_k_index[5965] = 27713;
mem_k_index[5966] = 27715;
mem_k_index[5967] = 27718;
mem_k_index[5968] = 27720;
mem_k_index[5969] = 27723;
mem_k_index[5970] = 27725;
mem_k_index[5971] = 27728;
mem_k_index[5972] = 27730;
mem_k_index[5973] = 27733;
mem_k_index[5974] = 27736;
mem_k_index[5975] = 27738;
mem_k_index[5976] = 27741;
mem_k_index[5977] = 27743;
mem_k_index[5978] = 27746;
mem_k_index[5979] = 27748;
mem_k_index[5980] = 27751;
mem_k_index[5981] = 27753;
mem_k_index[5982] = 27756;
mem_k_index[5983] = 27758;
mem_k_index[5984] = 27761;
mem_k_index[5985] = 27763;
mem_k_index[5986] = 27766;
mem_k_index[5987] = 27768;
mem_k_index[5988] = 27771;
mem_k_index[5989] = 27773;
mem_k_index[5990] = 27776;
mem_k_index[5991] = 27778;
mem_k_index[5992] = 27781;
mem_k_index[5993] = 27783;
mem_k_index[5994] = 27786;
mem_k_index[5995] = 27788;
mem_k_index[5996] = 27791;
mem_k_index[5997] = 27793;
mem_k_index[5998] = 27796;
mem_k_index[5999] = 27798;
mem_k_index[6000] = 27801;
mem_k_index[6001] = 27803;
mem_k_index[6002] = 27806;
mem_k_index[6003] = 27808;
mem_k_index[6004] = 27811;
mem_k_index[6005] = 27813;
mem_k_index[6006] = 27816;
mem_k_index[6007] = 27818;
mem_k_index[6008] = 27821;
mem_k_index[6009] = 27823;
mem_k_index[6010] = 27826;
mem_k_index[6011] = 27828;
mem_k_index[6012] = 27831;
mem_k_index[6013] = 27833;
mem_k_index[6014] = 27836;
mem_k_index[6015] = 27838;
mem_k_index[6016] = 28160;
mem_k_index[6017] = 28162;
mem_k_index[6018] = 28165;
mem_k_index[6019] = 28167;
mem_k_index[6020] = 28170;
mem_k_index[6021] = 28172;
mem_k_index[6022] = 28175;
mem_k_index[6023] = 28177;
mem_k_index[6024] = 28180;
mem_k_index[6025] = 28182;
mem_k_index[6026] = 28185;
mem_k_index[6027] = 28187;
mem_k_index[6028] = 28190;
mem_k_index[6029] = 28192;
mem_k_index[6030] = 28195;
mem_k_index[6031] = 28197;
mem_k_index[6032] = 28200;
mem_k_index[6033] = 28202;
mem_k_index[6034] = 28205;
mem_k_index[6035] = 28207;
mem_k_index[6036] = 28210;
mem_k_index[6037] = 28212;
mem_k_index[6038] = 28215;
mem_k_index[6039] = 28217;
mem_k_index[6040] = 28220;
mem_k_index[6041] = 28222;
mem_k_index[6042] = 28225;
mem_k_index[6043] = 28227;
mem_k_index[6044] = 28230;
mem_k_index[6045] = 28232;
mem_k_index[6046] = 28235;
mem_k_index[6047] = 28237;
mem_k_index[6048] = 28240;
mem_k_index[6049] = 28242;
mem_k_index[6050] = 28245;
mem_k_index[6051] = 28247;
mem_k_index[6052] = 28250;
mem_k_index[6053] = 28252;
mem_k_index[6054] = 28255;
mem_k_index[6055] = 28257;
mem_k_index[6056] = 28260;
mem_k_index[6057] = 28262;
mem_k_index[6058] = 28265;
mem_k_index[6059] = 28268;
mem_k_index[6060] = 28270;
mem_k_index[6061] = 28273;
mem_k_index[6062] = 28275;
mem_k_index[6063] = 28278;
mem_k_index[6064] = 28280;
mem_k_index[6065] = 28283;
mem_k_index[6066] = 28285;
mem_k_index[6067] = 28288;
mem_k_index[6068] = 28290;
mem_k_index[6069] = 28293;
mem_k_index[6070] = 28295;
mem_k_index[6071] = 28298;
mem_k_index[6072] = 28300;
mem_k_index[6073] = 28303;
mem_k_index[6074] = 28305;
mem_k_index[6075] = 28308;
mem_k_index[6076] = 28310;
mem_k_index[6077] = 28313;
mem_k_index[6078] = 28315;
mem_k_index[6079] = 28318;
mem_k_index[6080] = 28320;
mem_k_index[6081] = 28323;
mem_k_index[6082] = 28325;
mem_k_index[6083] = 28328;
mem_k_index[6084] = 28330;
mem_k_index[6085] = 28333;
mem_k_index[6086] = 28335;
mem_k_index[6087] = 28338;
mem_k_index[6088] = 28340;
mem_k_index[6089] = 28343;
mem_k_index[6090] = 28345;
mem_k_index[6091] = 28348;
mem_k_index[6092] = 28350;
mem_k_index[6093] = 28353;
mem_k_index[6094] = 28355;
mem_k_index[6095] = 28358;
mem_k_index[6096] = 28360;
mem_k_index[6097] = 28363;
mem_k_index[6098] = 28365;
mem_k_index[6099] = 28368;
mem_k_index[6100] = 28370;
mem_k_index[6101] = 28373;
mem_k_index[6102] = 28376;
mem_k_index[6103] = 28378;
mem_k_index[6104] = 28381;
mem_k_index[6105] = 28383;
mem_k_index[6106] = 28386;
mem_k_index[6107] = 28388;
mem_k_index[6108] = 28391;
mem_k_index[6109] = 28393;
mem_k_index[6110] = 28396;
mem_k_index[6111] = 28398;
mem_k_index[6112] = 28401;
mem_k_index[6113] = 28403;
mem_k_index[6114] = 28406;
mem_k_index[6115] = 28408;
mem_k_index[6116] = 28411;
mem_k_index[6117] = 28413;
mem_k_index[6118] = 28416;
mem_k_index[6119] = 28418;
mem_k_index[6120] = 28421;
mem_k_index[6121] = 28423;
mem_k_index[6122] = 28426;
mem_k_index[6123] = 28428;
mem_k_index[6124] = 28431;
mem_k_index[6125] = 28433;
mem_k_index[6126] = 28436;
mem_k_index[6127] = 28438;
mem_k_index[6128] = 28441;
mem_k_index[6129] = 28443;
mem_k_index[6130] = 28446;
mem_k_index[6131] = 28448;
mem_k_index[6132] = 28451;
mem_k_index[6133] = 28453;
mem_k_index[6134] = 28456;
mem_k_index[6135] = 28458;
mem_k_index[6136] = 28461;
mem_k_index[6137] = 28463;
mem_k_index[6138] = 28466;
mem_k_index[6139] = 28468;
mem_k_index[6140] = 28471;
mem_k_index[6141] = 28473;
mem_k_index[6142] = 28476;
mem_k_index[6143] = 28478;
mem_k_index[6144] = 28800;
mem_k_index[6145] = 28802;
mem_k_index[6146] = 28805;
mem_k_index[6147] = 28807;
mem_k_index[6148] = 28810;
mem_k_index[6149] = 28812;
mem_k_index[6150] = 28815;
mem_k_index[6151] = 28817;
mem_k_index[6152] = 28820;
mem_k_index[6153] = 28822;
mem_k_index[6154] = 28825;
mem_k_index[6155] = 28827;
mem_k_index[6156] = 28830;
mem_k_index[6157] = 28832;
mem_k_index[6158] = 28835;
mem_k_index[6159] = 28837;
mem_k_index[6160] = 28840;
mem_k_index[6161] = 28842;
mem_k_index[6162] = 28845;
mem_k_index[6163] = 28847;
mem_k_index[6164] = 28850;
mem_k_index[6165] = 28852;
mem_k_index[6166] = 28855;
mem_k_index[6167] = 28857;
mem_k_index[6168] = 28860;
mem_k_index[6169] = 28862;
mem_k_index[6170] = 28865;
mem_k_index[6171] = 28867;
mem_k_index[6172] = 28870;
mem_k_index[6173] = 28872;
mem_k_index[6174] = 28875;
mem_k_index[6175] = 28877;
mem_k_index[6176] = 28880;
mem_k_index[6177] = 28882;
mem_k_index[6178] = 28885;
mem_k_index[6179] = 28887;
mem_k_index[6180] = 28890;
mem_k_index[6181] = 28892;
mem_k_index[6182] = 28895;
mem_k_index[6183] = 28897;
mem_k_index[6184] = 28900;
mem_k_index[6185] = 28902;
mem_k_index[6186] = 28905;
mem_k_index[6187] = 28908;
mem_k_index[6188] = 28910;
mem_k_index[6189] = 28913;
mem_k_index[6190] = 28915;
mem_k_index[6191] = 28918;
mem_k_index[6192] = 28920;
mem_k_index[6193] = 28923;
mem_k_index[6194] = 28925;
mem_k_index[6195] = 28928;
mem_k_index[6196] = 28930;
mem_k_index[6197] = 28933;
mem_k_index[6198] = 28935;
mem_k_index[6199] = 28938;
mem_k_index[6200] = 28940;
mem_k_index[6201] = 28943;
mem_k_index[6202] = 28945;
mem_k_index[6203] = 28948;
mem_k_index[6204] = 28950;
mem_k_index[6205] = 28953;
mem_k_index[6206] = 28955;
mem_k_index[6207] = 28958;
mem_k_index[6208] = 28960;
mem_k_index[6209] = 28963;
mem_k_index[6210] = 28965;
mem_k_index[6211] = 28968;
mem_k_index[6212] = 28970;
mem_k_index[6213] = 28973;
mem_k_index[6214] = 28975;
mem_k_index[6215] = 28978;
mem_k_index[6216] = 28980;
mem_k_index[6217] = 28983;
mem_k_index[6218] = 28985;
mem_k_index[6219] = 28988;
mem_k_index[6220] = 28990;
mem_k_index[6221] = 28993;
mem_k_index[6222] = 28995;
mem_k_index[6223] = 28998;
mem_k_index[6224] = 29000;
mem_k_index[6225] = 29003;
mem_k_index[6226] = 29005;
mem_k_index[6227] = 29008;
mem_k_index[6228] = 29010;
mem_k_index[6229] = 29013;
mem_k_index[6230] = 29016;
mem_k_index[6231] = 29018;
mem_k_index[6232] = 29021;
mem_k_index[6233] = 29023;
mem_k_index[6234] = 29026;
mem_k_index[6235] = 29028;
mem_k_index[6236] = 29031;
mem_k_index[6237] = 29033;
mem_k_index[6238] = 29036;
mem_k_index[6239] = 29038;
mem_k_index[6240] = 29041;
mem_k_index[6241] = 29043;
mem_k_index[6242] = 29046;
mem_k_index[6243] = 29048;
mem_k_index[6244] = 29051;
mem_k_index[6245] = 29053;
mem_k_index[6246] = 29056;
mem_k_index[6247] = 29058;
mem_k_index[6248] = 29061;
mem_k_index[6249] = 29063;
mem_k_index[6250] = 29066;
mem_k_index[6251] = 29068;
mem_k_index[6252] = 29071;
mem_k_index[6253] = 29073;
mem_k_index[6254] = 29076;
mem_k_index[6255] = 29078;
mem_k_index[6256] = 29081;
mem_k_index[6257] = 29083;
mem_k_index[6258] = 29086;
mem_k_index[6259] = 29088;
mem_k_index[6260] = 29091;
mem_k_index[6261] = 29093;
mem_k_index[6262] = 29096;
mem_k_index[6263] = 29098;
mem_k_index[6264] = 29101;
mem_k_index[6265] = 29103;
mem_k_index[6266] = 29106;
mem_k_index[6267] = 29108;
mem_k_index[6268] = 29111;
mem_k_index[6269] = 29113;
mem_k_index[6270] = 29116;
mem_k_index[6271] = 29118;
mem_k_index[6272] = 29440;
mem_k_index[6273] = 29442;
mem_k_index[6274] = 29445;
mem_k_index[6275] = 29447;
mem_k_index[6276] = 29450;
mem_k_index[6277] = 29452;
mem_k_index[6278] = 29455;
mem_k_index[6279] = 29457;
mem_k_index[6280] = 29460;
mem_k_index[6281] = 29462;
mem_k_index[6282] = 29465;
mem_k_index[6283] = 29467;
mem_k_index[6284] = 29470;
mem_k_index[6285] = 29472;
mem_k_index[6286] = 29475;
mem_k_index[6287] = 29477;
mem_k_index[6288] = 29480;
mem_k_index[6289] = 29482;
mem_k_index[6290] = 29485;
mem_k_index[6291] = 29487;
mem_k_index[6292] = 29490;
mem_k_index[6293] = 29492;
mem_k_index[6294] = 29495;
mem_k_index[6295] = 29497;
mem_k_index[6296] = 29500;
mem_k_index[6297] = 29502;
mem_k_index[6298] = 29505;
mem_k_index[6299] = 29507;
mem_k_index[6300] = 29510;
mem_k_index[6301] = 29512;
mem_k_index[6302] = 29515;
mem_k_index[6303] = 29517;
mem_k_index[6304] = 29520;
mem_k_index[6305] = 29522;
mem_k_index[6306] = 29525;
mem_k_index[6307] = 29527;
mem_k_index[6308] = 29530;
mem_k_index[6309] = 29532;
mem_k_index[6310] = 29535;
mem_k_index[6311] = 29537;
mem_k_index[6312] = 29540;
mem_k_index[6313] = 29542;
mem_k_index[6314] = 29545;
mem_k_index[6315] = 29548;
mem_k_index[6316] = 29550;
mem_k_index[6317] = 29553;
mem_k_index[6318] = 29555;
mem_k_index[6319] = 29558;
mem_k_index[6320] = 29560;
mem_k_index[6321] = 29563;
mem_k_index[6322] = 29565;
mem_k_index[6323] = 29568;
mem_k_index[6324] = 29570;
mem_k_index[6325] = 29573;
mem_k_index[6326] = 29575;
mem_k_index[6327] = 29578;
mem_k_index[6328] = 29580;
mem_k_index[6329] = 29583;
mem_k_index[6330] = 29585;
mem_k_index[6331] = 29588;
mem_k_index[6332] = 29590;
mem_k_index[6333] = 29593;
mem_k_index[6334] = 29595;
mem_k_index[6335] = 29598;
mem_k_index[6336] = 29600;
mem_k_index[6337] = 29603;
mem_k_index[6338] = 29605;
mem_k_index[6339] = 29608;
mem_k_index[6340] = 29610;
mem_k_index[6341] = 29613;
mem_k_index[6342] = 29615;
mem_k_index[6343] = 29618;
mem_k_index[6344] = 29620;
mem_k_index[6345] = 29623;
mem_k_index[6346] = 29625;
mem_k_index[6347] = 29628;
mem_k_index[6348] = 29630;
mem_k_index[6349] = 29633;
mem_k_index[6350] = 29635;
mem_k_index[6351] = 29638;
mem_k_index[6352] = 29640;
mem_k_index[6353] = 29643;
mem_k_index[6354] = 29645;
mem_k_index[6355] = 29648;
mem_k_index[6356] = 29650;
mem_k_index[6357] = 29653;
mem_k_index[6358] = 29656;
mem_k_index[6359] = 29658;
mem_k_index[6360] = 29661;
mem_k_index[6361] = 29663;
mem_k_index[6362] = 29666;
mem_k_index[6363] = 29668;
mem_k_index[6364] = 29671;
mem_k_index[6365] = 29673;
mem_k_index[6366] = 29676;
mem_k_index[6367] = 29678;
mem_k_index[6368] = 29681;
mem_k_index[6369] = 29683;
mem_k_index[6370] = 29686;
mem_k_index[6371] = 29688;
mem_k_index[6372] = 29691;
mem_k_index[6373] = 29693;
mem_k_index[6374] = 29696;
mem_k_index[6375] = 29698;
mem_k_index[6376] = 29701;
mem_k_index[6377] = 29703;
mem_k_index[6378] = 29706;
mem_k_index[6379] = 29708;
mem_k_index[6380] = 29711;
mem_k_index[6381] = 29713;
mem_k_index[6382] = 29716;
mem_k_index[6383] = 29718;
mem_k_index[6384] = 29721;
mem_k_index[6385] = 29723;
mem_k_index[6386] = 29726;
mem_k_index[6387] = 29728;
mem_k_index[6388] = 29731;
mem_k_index[6389] = 29733;
mem_k_index[6390] = 29736;
mem_k_index[6391] = 29738;
mem_k_index[6392] = 29741;
mem_k_index[6393] = 29743;
mem_k_index[6394] = 29746;
mem_k_index[6395] = 29748;
mem_k_index[6396] = 29751;
mem_k_index[6397] = 29753;
mem_k_index[6398] = 29756;
mem_k_index[6399] = 29758;
mem_k_index[6400] = 30080;
mem_k_index[6401] = 30082;
mem_k_index[6402] = 30085;
mem_k_index[6403] = 30087;
mem_k_index[6404] = 30090;
mem_k_index[6405] = 30092;
mem_k_index[6406] = 30095;
mem_k_index[6407] = 30097;
mem_k_index[6408] = 30100;
mem_k_index[6409] = 30102;
mem_k_index[6410] = 30105;
mem_k_index[6411] = 30107;
mem_k_index[6412] = 30110;
mem_k_index[6413] = 30112;
mem_k_index[6414] = 30115;
mem_k_index[6415] = 30117;
mem_k_index[6416] = 30120;
mem_k_index[6417] = 30122;
mem_k_index[6418] = 30125;
mem_k_index[6419] = 30127;
mem_k_index[6420] = 30130;
mem_k_index[6421] = 30132;
mem_k_index[6422] = 30135;
mem_k_index[6423] = 30137;
mem_k_index[6424] = 30140;
mem_k_index[6425] = 30142;
mem_k_index[6426] = 30145;
mem_k_index[6427] = 30147;
mem_k_index[6428] = 30150;
mem_k_index[6429] = 30152;
mem_k_index[6430] = 30155;
mem_k_index[6431] = 30157;
mem_k_index[6432] = 30160;
mem_k_index[6433] = 30162;
mem_k_index[6434] = 30165;
mem_k_index[6435] = 30167;
mem_k_index[6436] = 30170;
mem_k_index[6437] = 30172;
mem_k_index[6438] = 30175;
mem_k_index[6439] = 30177;
mem_k_index[6440] = 30180;
mem_k_index[6441] = 30182;
mem_k_index[6442] = 30185;
mem_k_index[6443] = 30188;
mem_k_index[6444] = 30190;
mem_k_index[6445] = 30193;
mem_k_index[6446] = 30195;
mem_k_index[6447] = 30198;
mem_k_index[6448] = 30200;
mem_k_index[6449] = 30203;
mem_k_index[6450] = 30205;
mem_k_index[6451] = 30208;
mem_k_index[6452] = 30210;
mem_k_index[6453] = 30213;
mem_k_index[6454] = 30215;
mem_k_index[6455] = 30218;
mem_k_index[6456] = 30220;
mem_k_index[6457] = 30223;
mem_k_index[6458] = 30225;
mem_k_index[6459] = 30228;
mem_k_index[6460] = 30230;
mem_k_index[6461] = 30233;
mem_k_index[6462] = 30235;
mem_k_index[6463] = 30238;
mem_k_index[6464] = 30240;
mem_k_index[6465] = 30243;
mem_k_index[6466] = 30245;
mem_k_index[6467] = 30248;
mem_k_index[6468] = 30250;
mem_k_index[6469] = 30253;
mem_k_index[6470] = 30255;
mem_k_index[6471] = 30258;
mem_k_index[6472] = 30260;
mem_k_index[6473] = 30263;
mem_k_index[6474] = 30265;
mem_k_index[6475] = 30268;
mem_k_index[6476] = 30270;
mem_k_index[6477] = 30273;
mem_k_index[6478] = 30275;
mem_k_index[6479] = 30278;
mem_k_index[6480] = 30280;
mem_k_index[6481] = 30283;
mem_k_index[6482] = 30285;
mem_k_index[6483] = 30288;
mem_k_index[6484] = 30290;
mem_k_index[6485] = 30293;
mem_k_index[6486] = 30296;
mem_k_index[6487] = 30298;
mem_k_index[6488] = 30301;
mem_k_index[6489] = 30303;
mem_k_index[6490] = 30306;
mem_k_index[6491] = 30308;
mem_k_index[6492] = 30311;
mem_k_index[6493] = 30313;
mem_k_index[6494] = 30316;
mem_k_index[6495] = 30318;
mem_k_index[6496] = 30321;
mem_k_index[6497] = 30323;
mem_k_index[6498] = 30326;
mem_k_index[6499] = 30328;
mem_k_index[6500] = 30331;
mem_k_index[6501] = 30333;
mem_k_index[6502] = 30336;
mem_k_index[6503] = 30338;
mem_k_index[6504] = 30341;
mem_k_index[6505] = 30343;
mem_k_index[6506] = 30346;
mem_k_index[6507] = 30348;
mem_k_index[6508] = 30351;
mem_k_index[6509] = 30353;
mem_k_index[6510] = 30356;
mem_k_index[6511] = 30358;
mem_k_index[6512] = 30361;
mem_k_index[6513] = 30363;
mem_k_index[6514] = 30366;
mem_k_index[6515] = 30368;
mem_k_index[6516] = 30371;
mem_k_index[6517] = 30373;
mem_k_index[6518] = 30376;
mem_k_index[6519] = 30378;
mem_k_index[6520] = 30381;
mem_k_index[6521] = 30383;
mem_k_index[6522] = 30386;
mem_k_index[6523] = 30388;
mem_k_index[6524] = 30391;
mem_k_index[6525] = 30393;
mem_k_index[6526] = 30396;
mem_k_index[6527] = 30398;
mem_k_index[6528] = 30400;
mem_k_index[6529] = 30402;
mem_k_index[6530] = 30405;
mem_k_index[6531] = 30407;
mem_k_index[6532] = 30410;
mem_k_index[6533] = 30412;
mem_k_index[6534] = 30415;
mem_k_index[6535] = 30417;
mem_k_index[6536] = 30420;
mem_k_index[6537] = 30422;
mem_k_index[6538] = 30425;
mem_k_index[6539] = 30427;
mem_k_index[6540] = 30430;
mem_k_index[6541] = 30432;
mem_k_index[6542] = 30435;
mem_k_index[6543] = 30437;
mem_k_index[6544] = 30440;
mem_k_index[6545] = 30442;
mem_k_index[6546] = 30445;
mem_k_index[6547] = 30447;
mem_k_index[6548] = 30450;
mem_k_index[6549] = 30452;
mem_k_index[6550] = 30455;
mem_k_index[6551] = 30457;
mem_k_index[6552] = 30460;
mem_k_index[6553] = 30462;
mem_k_index[6554] = 30465;
mem_k_index[6555] = 30467;
mem_k_index[6556] = 30470;
mem_k_index[6557] = 30472;
mem_k_index[6558] = 30475;
mem_k_index[6559] = 30477;
mem_k_index[6560] = 30480;
mem_k_index[6561] = 30482;
mem_k_index[6562] = 30485;
mem_k_index[6563] = 30487;
mem_k_index[6564] = 30490;
mem_k_index[6565] = 30492;
mem_k_index[6566] = 30495;
mem_k_index[6567] = 30497;
mem_k_index[6568] = 30500;
mem_k_index[6569] = 30502;
mem_k_index[6570] = 30505;
mem_k_index[6571] = 30508;
mem_k_index[6572] = 30510;
mem_k_index[6573] = 30513;
mem_k_index[6574] = 30515;
mem_k_index[6575] = 30518;
mem_k_index[6576] = 30520;
mem_k_index[6577] = 30523;
mem_k_index[6578] = 30525;
mem_k_index[6579] = 30528;
mem_k_index[6580] = 30530;
mem_k_index[6581] = 30533;
mem_k_index[6582] = 30535;
mem_k_index[6583] = 30538;
mem_k_index[6584] = 30540;
mem_k_index[6585] = 30543;
mem_k_index[6586] = 30545;
mem_k_index[6587] = 30548;
mem_k_index[6588] = 30550;
mem_k_index[6589] = 30553;
mem_k_index[6590] = 30555;
mem_k_index[6591] = 30558;
mem_k_index[6592] = 30560;
mem_k_index[6593] = 30563;
mem_k_index[6594] = 30565;
mem_k_index[6595] = 30568;
mem_k_index[6596] = 30570;
mem_k_index[6597] = 30573;
mem_k_index[6598] = 30575;
mem_k_index[6599] = 30578;
mem_k_index[6600] = 30580;
mem_k_index[6601] = 30583;
mem_k_index[6602] = 30585;
mem_k_index[6603] = 30588;
mem_k_index[6604] = 30590;
mem_k_index[6605] = 30593;
mem_k_index[6606] = 30595;
mem_k_index[6607] = 30598;
mem_k_index[6608] = 30600;
mem_k_index[6609] = 30603;
mem_k_index[6610] = 30605;
mem_k_index[6611] = 30608;
mem_k_index[6612] = 30610;
mem_k_index[6613] = 30613;
mem_k_index[6614] = 30616;
mem_k_index[6615] = 30618;
mem_k_index[6616] = 30621;
mem_k_index[6617] = 30623;
mem_k_index[6618] = 30626;
mem_k_index[6619] = 30628;
mem_k_index[6620] = 30631;
mem_k_index[6621] = 30633;
mem_k_index[6622] = 30636;
mem_k_index[6623] = 30638;
mem_k_index[6624] = 30641;
mem_k_index[6625] = 30643;
mem_k_index[6626] = 30646;
mem_k_index[6627] = 30648;
mem_k_index[6628] = 30651;
mem_k_index[6629] = 30653;
mem_k_index[6630] = 30656;
mem_k_index[6631] = 30658;
mem_k_index[6632] = 30661;
mem_k_index[6633] = 30663;
mem_k_index[6634] = 30666;
mem_k_index[6635] = 30668;
mem_k_index[6636] = 30671;
mem_k_index[6637] = 30673;
mem_k_index[6638] = 30676;
mem_k_index[6639] = 30678;
mem_k_index[6640] = 30681;
mem_k_index[6641] = 30683;
mem_k_index[6642] = 30686;
mem_k_index[6643] = 30688;
mem_k_index[6644] = 30691;
mem_k_index[6645] = 30693;
mem_k_index[6646] = 30696;
mem_k_index[6647] = 30698;
mem_k_index[6648] = 30701;
mem_k_index[6649] = 30703;
mem_k_index[6650] = 30706;
mem_k_index[6651] = 30708;
mem_k_index[6652] = 30711;
mem_k_index[6653] = 30713;
mem_k_index[6654] = 30716;
mem_k_index[6655] = 30718;
mem_k_index[6656] = 31040;
mem_k_index[6657] = 31042;
mem_k_index[6658] = 31045;
mem_k_index[6659] = 31047;
mem_k_index[6660] = 31050;
mem_k_index[6661] = 31052;
mem_k_index[6662] = 31055;
mem_k_index[6663] = 31057;
mem_k_index[6664] = 31060;
mem_k_index[6665] = 31062;
mem_k_index[6666] = 31065;
mem_k_index[6667] = 31067;
mem_k_index[6668] = 31070;
mem_k_index[6669] = 31072;
mem_k_index[6670] = 31075;
mem_k_index[6671] = 31077;
mem_k_index[6672] = 31080;
mem_k_index[6673] = 31082;
mem_k_index[6674] = 31085;
mem_k_index[6675] = 31087;
mem_k_index[6676] = 31090;
mem_k_index[6677] = 31092;
mem_k_index[6678] = 31095;
mem_k_index[6679] = 31097;
mem_k_index[6680] = 31100;
mem_k_index[6681] = 31102;
mem_k_index[6682] = 31105;
mem_k_index[6683] = 31107;
mem_k_index[6684] = 31110;
mem_k_index[6685] = 31112;
mem_k_index[6686] = 31115;
mem_k_index[6687] = 31117;
mem_k_index[6688] = 31120;
mem_k_index[6689] = 31122;
mem_k_index[6690] = 31125;
mem_k_index[6691] = 31127;
mem_k_index[6692] = 31130;
mem_k_index[6693] = 31132;
mem_k_index[6694] = 31135;
mem_k_index[6695] = 31137;
mem_k_index[6696] = 31140;
mem_k_index[6697] = 31142;
mem_k_index[6698] = 31145;
mem_k_index[6699] = 31148;
mem_k_index[6700] = 31150;
mem_k_index[6701] = 31153;
mem_k_index[6702] = 31155;
mem_k_index[6703] = 31158;
mem_k_index[6704] = 31160;
mem_k_index[6705] = 31163;
mem_k_index[6706] = 31165;
mem_k_index[6707] = 31168;
mem_k_index[6708] = 31170;
mem_k_index[6709] = 31173;
mem_k_index[6710] = 31175;
mem_k_index[6711] = 31178;
mem_k_index[6712] = 31180;
mem_k_index[6713] = 31183;
mem_k_index[6714] = 31185;
mem_k_index[6715] = 31188;
mem_k_index[6716] = 31190;
mem_k_index[6717] = 31193;
mem_k_index[6718] = 31195;
mem_k_index[6719] = 31198;
mem_k_index[6720] = 31200;
mem_k_index[6721] = 31203;
mem_k_index[6722] = 31205;
mem_k_index[6723] = 31208;
mem_k_index[6724] = 31210;
mem_k_index[6725] = 31213;
mem_k_index[6726] = 31215;
mem_k_index[6727] = 31218;
mem_k_index[6728] = 31220;
mem_k_index[6729] = 31223;
mem_k_index[6730] = 31225;
mem_k_index[6731] = 31228;
mem_k_index[6732] = 31230;
mem_k_index[6733] = 31233;
mem_k_index[6734] = 31235;
mem_k_index[6735] = 31238;
mem_k_index[6736] = 31240;
mem_k_index[6737] = 31243;
mem_k_index[6738] = 31245;
mem_k_index[6739] = 31248;
mem_k_index[6740] = 31250;
mem_k_index[6741] = 31253;
mem_k_index[6742] = 31256;
mem_k_index[6743] = 31258;
mem_k_index[6744] = 31261;
mem_k_index[6745] = 31263;
mem_k_index[6746] = 31266;
mem_k_index[6747] = 31268;
mem_k_index[6748] = 31271;
mem_k_index[6749] = 31273;
mem_k_index[6750] = 31276;
mem_k_index[6751] = 31278;
mem_k_index[6752] = 31281;
mem_k_index[6753] = 31283;
mem_k_index[6754] = 31286;
mem_k_index[6755] = 31288;
mem_k_index[6756] = 31291;
mem_k_index[6757] = 31293;
mem_k_index[6758] = 31296;
mem_k_index[6759] = 31298;
mem_k_index[6760] = 31301;
mem_k_index[6761] = 31303;
mem_k_index[6762] = 31306;
mem_k_index[6763] = 31308;
mem_k_index[6764] = 31311;
mem_k_index[6765] = 31313;
mem_k_index[6766] = 31316;
mem_k_index[6767] = 31318;
mem_k_index[6768] = 31321;
mem_k_index[6769] = 31323;
mem_k_index[6770] = 31326;
mem_k_index[6771] = 31328;
mem_k_index[6772] = 31331;
mem_k_index[6773] = 31333;
mem_k_index[6774] = 31336;
mem_k_index[6775] = 31338;
mem_k_index[6776] = 31341;
mem_k_index[6777] = 31343;
mem_k_index[6778] = 31346;
mem_k_index[6779] = 31348;
mem_k_index[6780] = 31351;
mem_k_index[6781] = 31353;
mem_k_index[6782] = 31356;
mem_k_index[6783] = 31358;
mem_k_index[6784] = 31680;
mem_k_index[6785] = 31682;
mem_k_index[6786] = 31685;
mem_k_index[6787] = 31687;
mem_k_index[6788] = 31690;
mem_k_index[6789] = 31692;
mem_k_index[6790] = 31695;
mem_k_index[6791] = 31697;
mem_k_index[6792] = 31700;
mem_k_index[6793] = 31702;
mem_k_index[6794] = 31705;
mem_k_index[6795] = 31707;
mem_k_index[6796] = 31710;
mem_k_index[6797] = 31712;
mem_k_index[6798] = 31715;
mem_k_index[6799] = 31717;
mem_k_index[6800] = 31720;
mem_k_index[6801] = 31722;
mem_k_index[6802] = 31725;
mem_k_index[6803] = 31727;
mem_k_index[6804] = 31730;
mem_k_index[6805] = 31732;
mem_k_index[6806] = 31735;
mem_k_index[6807] = 31737;
mem_k_index[6808] = 31740;
mem_k_index[6809] = 31742;
mem_k_index[6810] = 31745;
mem_k_index[6811] = 31747;
mem_k_index[6812] = 31750;
mem_k_index[6813] = 31752;
mem_k_index[6814] = 31755;
mem_k_index[6815] = 31757;
mem_k_index[6816] = 31760;
mem_k_index[6817] = 31762;
mem_k_index[6818] = 31765;
mem_k_index[6819] = 31767;
mem_k_index[6820] = 31770;
mem_k_index[6821] = 31772;
mem_k_index[6822] = 31775;
mem_k_index[6823] = 31777;
mem_k_index[6824] = 31780;
mem_k_index[6825] = 31782;
mem_k_index[6826] = 31785;
mem_k_index[6827] = 31788;
mem_k_index[6828] = 31790;
mem_k_index[6829] = 31793;
mem_k_index[6830] = 31795;
mem_k_index[6831] = 31798;
mem_k_index[6832] = 31800;
mem_k_index[6833] = 31803;
mem_k_index[6834] = 31805;
mem_k_index[6835] = 31808;
mem_k_index[6836] = 31810;
mem_k_index[6837] = 31813;
mem_k_index[6838] = 31815;
mem_k_index[6839] = 31818;
mem_k_index[6840] = 31820;
mem_k_index[6841] = 31823;
mem_k_index[6842] = 31825;
mem_k_index[6843] = 31828;
mem_k_index[6844] = 31830;
mem_k_index[6845] = 31833;
mem_k_index[6846] = 31835;
mem_k_index[6847] = 31838;
mem_k_index[6848] = 31840;
mem_k_index[6849] = 31843;
mem_k_index[6850] = 31845;
mem_k_index[6851] = 31848;
mem_k_index[6852] = 31850;
mem_k_index[6853] = 31853;
mem_k_index[6854] = 31855;
mem_k_index[6855] = 31858;
mem_k_index[6856] = 31860;
mem_k_index[6857] = 31863;
mem_k_index[6858] = 31865;
mem_k_index[6859] = 31868;
mem_k_index[6860] = 31870;
mem_k_index[6861] = 31873;
mem_k_index[6862] = 31875;
mem_k_index[6863] = 31878;
mem_k_index[6864] = 31880;
mem_k_index[6865] = 31883;
mem_k_index[6866] = 31885;
mem_k_index[6867] = 31888;
mem_k_index[6868] = 31890;
mem_k_index[6869] = 31893;
mem_k_index[6870] = 31896;
mem_k_index[6871] = 31898;
mem_k_index[6872] = 31901;
mem_k_index[6873] = 31903;
mem_k_index[6874] = 31906;
mem_k_index[6875] = 31908;
mem_k_index[6876] = 31911;
mem_k_index[6877] = 31913;
mem_k_index[6878] = 31916;
mem_k_index[6879] = 31918;
mem_k_index[6880] = 31921;
mem_k_index[6881] = 31923;
mem_k_index[6882] = 31926;
mem_k_index[6883] = 31928;
mem_k_index[6884] = 31931;
mem_k_index[6885] = 31933;
mem_k_index[6886] = 31936;
mem_k_index[6887] = 31938;
mem_k_index[6888] = 31941;
mem_k_index[6889] = 31943;
mem_k_index[6890] = 31946;
mem_k_index[6891] = 31948;
mem_k_index[6892] = 31951;
mem_k_index[6893] = 31953;
mem_k_index[6894] = 31956;
mem_k_index[6895] = 31958;
mem_k_index[6896] = 31961;
mem_k_index[6897] = 31963;
mem_k_index[6898] = 31966;
mem_k_index[6899] = 31968;
mem_k_index[6900] = 31971;
mem_k_index[6901] = 31973;
mem_k_index[6902] = 31976;
mem_k_index[6903] = 31978;
mem_k_index[6904] = 31981;
mem_k_index[6905] = 31983;
mem_k_index[6906] = 31986;
mem_k_index[6907] = 31988;
mem_k_index[6908] = 31991;
mem_k_index[6909] = 31993;
mem_k_index[6910] = 31996;
mem_k_index[6911] = 31998;
mem_k_index[6912] = 32320;
mem_k_index[6913] = 32322;
mem_k_index[6914] = 32325;
mem_k_index[6915] = 32327;
mem_k_index[6916] = 32330;
mem_k_index[6917] = 32332;
mem_k_index[6918] = 32335;
mem_k_index[6919] = 32337;
mem_k_index[6920] = 32340;
mem_k_index[6921] = 32342;
mem_k_index[6922] = 32345;
mem_k_index[6923] = 32347;
mem_k_index[6924] = 32350;
mem_k_index[6925] = 32352;
mem_k_index[6926] = 32355;
mem_k_index[6927] = 32357;
mem_k_index[6928] = 32360;
mem_k_index[6929] = 32362;
mem_k_index[6930] = 32365;
mem_k_index[6931] = 32367;
mem_k_index[6932] = 32370;
mem_k_index[6933] = 32372;
mem_k_index[6934] = 32375;
mem_k_index[6935] = 32377;
mem_k_index[6936] = 32380;
mem_k_index[6937] = 32382;
mem_k_index[6938] = 32385;
mem_k_index[6939] = 32387;
mem_k_index[6940] = 32390;
mem_k_index[6941] = 32392;
mem_k_index[6942] = 32395;
mem_k_index[6943] = 32397;
mem_k_index[6944] = 32400;
mem_k_index[6945] = 32402;
mem_k_index[6946] = 32405;
mem_k_index[6947] = 32407;
mem_k_index[6948] = 32410;
mem_k_index[6949] = 32412;
mem_k_index[6950] = 32415;
mem_k_index[6951] = 32417;
mem_k_index[6952] = 32420;
mem_k_index[6953] = 32422;
mem_k_index[6954] = 32425;
mem_k_index[6955] = 32428;
mem_k_index[6956] = 32430;
mem_k_index[6957] = 32433;
mem_k_index[6958] = 32435;
mem_k_index[6959] = 32438;
mem_k_index[6960] = 32440;
mem_k_index[6961] = 32443;
mem_k_index[6962] = 32445;
mem_k_index[6963] = 32448;
mem_k_index[6964] = 32450;
mem_k_index[6965] = 32453;
mem_k_index[6966] = 32455;
mem_k_index[6967] = 32458;
mem_k_index[6968] = 32460;
mem_k_index[6969] = 32463;
mem_k_index[6970] = 32465;
mem_k_index[6971] = 32468;
mem_k_index[6972] = 32470;
mem_k_index[6973] = 32473;
mem_k_index[6974] = 32475;
mem_k_index[6975] = 32478;
mem_k_index[6976] = 32480;
mem_k_index[6977] = 32483;
mem_k_index[6978] = 32485;
mem_k_index[6979] = 32488;
mem_k_index[6980] = 32490;
mem_k_index[6981] = 32493;
mem_k_index[6982] = 32495;
mem_k_index[6983] = 32498;
mem_k_index[6984] = 32500;
mem_k_index[6985] = 32503;
mem_k_index[6986] = 32505;
mem_k_index[6987] = 32508;
mem_k_index[6988] = 32510;
mem_k_index[6989] = 32513;
mem_k_index[6990] = 32515;
mem_k_index[6991] = 32518;
mem_k_index[6992] = 32520;
mem_k_index[6993] = 32523;
mem_k_index[6994] = 32525;
mem_k_index[6995] = 32528;
mem_k_index[6996] = 32530;
mem_k_index[6997] = 32533;
mem_k_index[6998] = 32536;
mem_k_index[6999] = 32538;
mem_k_index[7000] = 32541;
mem_k_index[7001] = 32543;
mem_k_index[7002] = 32546;
mem_k_index[7003] = 32548;
mem_k_index[7004] = 32551;
mem_k_index[7005] = 32553;
mem_k_index[7006] = 32556;
mem_k_index[7007] = 32558;
mem_k_index[7008] = 32561;
mem_k_index[7009] = 32563;
mem_k_index[7010] = 32566;
mem_k_index[7011] = 32568;
mem_k_index[7012] = 32571;
mem_k_index[7013] = 32573;
mem_k_index[7014] = 32576;
mem_k_index[7015] = 32578;
mem_k_index[7016] = 32581;
mem_k_index[7017] = 32583;
mem_k_index[7018] = 32586;
mem_k_index[7019] = 32588;
mem_k_index[7020] = 32591;
mem_k_index[7021] = 32593;
mem_k_index[7022] = 32596;
mem_k_index[7023] = 32598;
mem_k_index[7024] = 32601;
mem_k_index[7025] = 32603;
mem_k_index[7026] = 32606;
mem_k_index[7027] = 32608;
mem_k_index[7028] = 32611;
mem_k_index[7029] = 32613;
mem_k_index[7030] = 32616;
mem_k_index[7031] = 32618;
mem_k_index[7032] = 32621;
mem_k_index[7033] = 32623;
mem_k_index[7034] = 32626;
mem_k_index[7035] = 32628;
mem_k_index[7036] = 32631;
mem_k_index[7037] = 32633;
mem_k_index[7038] = 32636;
mem_k_index[7039] = 32638;
mem_k_index[7040] = 32960;
mem_k_index[7041] = 32962;
mem_k_index[7042] = 32965;
mem_k_index[7043] = 32967;
mem_k_index[7044] = 32970;
mem_k_index[7045] = 32972;
mem_k_index[7046] = 32975;
mem_k_index[7047] = 32977;
mem_k_index[7048] = 32980;
mem_k_index[7049] = 32982;
mem_k_index[7050] = 32985;
mem_k_index[7051] = 32987;
mem_k_index[7052] = 32990;
mem_k_index[7053] = 32992;
mem_k_index[7054] = 32995;
mem_k_index[7055] = 32997;
mem_k_index[7056] = 33000;
mem_k_index[7057] = 33002;
mem_k_index[7058] = 33005;
mem_k_index[7059] = 33007;
mem_k_index[7060] = 33010;
mem_k_index[7061] = 33012;
mem_k_index[7062] = 33015;
mem_k_index[7063] = 33017;
mem_k_index[7064] = 33020;
mem_k_index[7065] = 33022;
mem_k_index[7066] = 33025;
mem_k_index[7067] = 33027;
mem_k_index[7068] = 33030;
mem_k_index[7069] = 33032;
mem_k_index[7070] = 33035;
mem_k_index[7071] = 33037;
mem_k_index[7072] = 33040;
mem_k_index[7073] = 33042;
mem_k_index[7074] = 33045;
mem_k_index[7075] = 33047;
mem_k_index[7076] = 33050;
mem_k_index[7077] = 33052;
mem_k_index[7078] = 33055;
mem_k_index[7079] = 33057;
mem_k_index[7080] = 33060;
mem_k_index[7081] = 33062;
mem_k_index[7082] = 33065;
mem_k_index[7083] = 33068;
mem_k_index[7084] = 33070;
mem_k_index[7085] = 33073;
mem_k_index[7086] = 33075;
mem_k_index[7087] = 33078;
mem_k_index[7088] = 33080;
mem_k_index[7089] = 33083;
mem_k_index[7090] = 33085;
mem_k_index[7091] = 33088;
mem_k_index[7092] = 33090;
mem_k_index[7093] = 33093;
mem_k_index[7094] = 33095;
mem_k_index[7095] = 33098;
mem_k_index[7096] = 33100;
mem_k_index[7097] = 33103;
mem_k_index[7098] = 33105;
mem_k_index[7099] = 33108;
mem_k_index[7100] = 33110;
mem_k_index[7101] = 33113;
mem_k_index[7102] = 33115;
mem_k_index[7103] = 33118;
mem_k_index[7104] = 33120;
mem_k_index[7105] = 33123;
mem_k_index[7106] = 33125;
mem_k_index[7107] = 33128;
mem_k_index[7108] = 33130;
mem_k_index[7109] = 33133;
mem_k_index[7110] = 33135;
mem_k_index[7111] = 33138;
mem_k_index[7112] = 33140;
mem_k_index[7113] = 33143;
mem_k_index[7114] = 33145;
mem_k_index[7115] = 33148;
mem_k_index[7116] = 33150;
mem_k_index[7117] = 33153;
mem_k_index[7118] = 33155;
mem_k_index[7119] = 33158;
mem_k_index[7120] = 33160;
mem_k_index[7121] = 33163;
mem_k_index[7122] = 33165;
mem_k_index[7123] = 33168;
mem_k_index[7124] = 33170;
mem_k_index[7125] = 33173;
mem_k_index[7126] = 33176;
mem_k_index[7127] = 33178;
mem_k_index[7128] = 33181;
mem_k_index[7129] = 33183;
mem_k_index[7130] = 33186;
mem_k_index[7131] = 33188;
mem_k_index[7132] = 33191;
mem_k_index[7133] = 33193;
mem_k_index[7134] = 33196;
mem_k_index[7135] = 33198;
mem_k_index[7136] = 33201;
mem_k_index[7137] = 33203;
mem_k_index[7138] = 33206;
mem_k_index[7139] = 33208;
mem_k_index[7140] = 33211;
mem_k_index[7141] = 33213;
mem_k_index[7142] = 33216;
mem_k_index[7143] = 33218;
mem_k_index[7144] = 33221;
mem_k_index[7145] = 33223;
mem_k_index[7146] = 33226;
mem_k_index[7147] = 33228;
mem_k_index[7148] = 33231;
mem_k_index[7149] = 33233;
mem_k_index[7150] = 33236;
mem_k_index[7151] = 33238;
mem_k_index[7152] = 33241;
mem_k_index[7153] = 33243;
mem_k_index[7154] = 33246;
mem_k_index[7155] = 33248;
mem_k_index[7156] = 33251;
mem_k_index[7157] = 33253;
mem_k_index[7158] = 33256;
mem_k_index[7159] = 33258;
mem_k_index[7160] = 33261;
mem_k_index[7161] = 33263;
mem_k_index[7162] = 33266;
mem_k_index[7163] = 33268;
mem_k_index[7164] = 33271;
mem_k_index[7165] = 33273;
mem_k_index[7166] = 33276;
mem_k_index[7167] = 33278;
mem_k_index[7168] = 33600;
mem_k_index[7169] = 33602;
mem_k_index[7170] = 33605;
mem_k_index[7171] = 33607;
mem_k_index[7172] = 33610;
mem_k_index[7173] = 33612;
mem_k_index[7174] = 33615;
mem_k_index[7175] = 33617;
mem_k_index[7176] = 33620;
mem_k_index[7177] = 33622;
mem_k_index[7178] = 33625;
mem_k_index[7179] = 33627;
mem_k_index[7180] = 33630;
mem_k_index[7181] = 33632;
mem_k_index[7182] = 33635;
mem_k_index[7183] = 33637;
mem_k_index[7184] = 33640;
mem_k_index[7185] = 33642;
mem_k_index[7186] = 33645;
mem_k_index[7187] = 33647;
mem_k_index[7188] = 33650;
mem_k_index[7189] = 33652;
mem_k_index[7190] = 33655;
mem_k_index[7191] = 33657;
mem_k_index[7192] = 33660;
mem_k_index[7193] = 33662;
mem_k_index[7194] = 33665;
mem_k_index[7195] = 33667;
mem_k_index[7196] = 33670;
mem_k_index[7197] = 33672;
mem_k_index[7198] = 33675;
mem_k_index[7199] = 33677;
mem_k_index[7200] = 33680;
mem_k_index[7201] = 33682;
mem_k_index[7202] = 33685;
mem_k_index[7203] = 33687;
mem_k_index[7204] = 33690;
mem_k_index[7205] = 33692;
mem_k_index[7206] = 33695;
mem_k_index[7207] = 33697;
mem_k_index[7208] = 33700;
mem_k_index[7209] = 33702;
mem_k_index[7210] = 33705;
mem_k_index[7211] = 33708;
mem_k_index[7212] = 33710;
mem_k_index[7213] = 33713;
mem_k_index[7214] = 33715;
mem_k_index[7215] = 33718;
mem_k_index[7216] = 33720;
mem_k_index[7217] = 33723;
mem_k_index[7218] = 33725;
mem_k_index[7219] = 33728;
mem_k_index[7220] = 33730;
mem_k_index[7221] = 33733;
mem_k_index[7222] = 33735;
mem_k_index[7223] = 33738;
mem_k_index[7224] = 33740;
mem_k_index[7225] = 33743;
mem_k_index[7226] = 33745;
mem_k_index[7227] = 33748;
mem_k_index[7228] = 33750;
mem_k_index[7229] = 33753;
mem_k_index[7230] = 33755;
mem_k_index[7231] = 33758;
mem_k_index[7232] = 33760;
mem_k_index[7233] = 33763;
mem_k_index[7234] = 33765;
mem_k_index[7235] = 33768;
mem_k_index[7236] = 33770;
mem_k_index[7237] = 33773;
mem_k_index[7238] = 33775;
mem_k_index[7239] = 33778;
mem_k_index[7240] = 33780;
mem_k_index[7241] = 33783;
mem_k_index[7242] = 33785;
mem_k_index[7243] = 33788;
mem_k_index[7244] = 33790;
mem_k_index[7245] = 33793;
mem_k_index[7246] = 33795;
mem_k_index[7247] = 33798;
mem_k_index[7248] = 33800;
mem_k_index[7249] = 33803;
mem_k_index[7250] = 33805;
mem_k_index[7251] = 33808;
mem_k_index[7252] = 33810;
mem_k_index[7253] = 33813;
mem_k_index[7254] = 33816;
mem_k_index[7255] = 33818;
mem_k_index[7256] = 33821;
mem_k_index[7257] = 33823;
mem_k_index[7258] = 33826;
mem_k_index[7259] = 33828;
mem_k_index[7260] = 33831;
mem_k_index[7261] = 33833;
mem_k_index[7262] = 33836;
mem_k_index[7263] = 33838;
mem_k_index[7264] = 33841;
mem_k_index[7265] = 33843;
mem_k_index[7266] = 33846;
mem_k_index[7267] = 33848;
mem_k_index[7268] = 33851;
mem_k_index[7269] = 33853;
mem_k_index[7270] = 33856;
mem_k_index[7271] = 33858;
mem_k_index[7272] = 33861;
mem_k_index[7273] = 33863;
mem_k_index[7274] = 33866;
mem_k_index[7275] = 33868;
mem_k_index[7276] = 33871;
mem_k_index[7277] = 33873;
mem_k_index[7278] = 33876;
mem_k_index[7279] = 33878;
mem_k_index[7280] = 33881;
mem_k_index[7281] = 33883;
mem_k_index[7282] = 33886;
mem_k_index[7283] = 33888;
mem_k_index[7284] = 33891;
mem_k_index[7285] = 33893;
mem_k_index[7286] = 33896;
mem_k_index[7287] = 33898;
mem_k_index[7288] = 33901;
mem_k_index[7289] = 33903;
mem_k_index[7290] = 33906;
mem_k_index[7291] = 33908;
mem_k_index[7292] = 33911;
mem_k_index[7293] = 33913;
mem_k_index[7294] = 33916;
mem_k_index[7295] = 33918;
mem_k_index[7296] = 34240;
mem_k_index[7297] = 34242;
mem_k_index[7298] = 34245;
mem_k_index[7299] = 34247;
mem_k_index[7300] = 34250;
mem_k_index[7301] = 34252;
mem_k_index[7302] = 34255;
mem_k_index[7303] = 34257;
mem_k_index[7304] = 34260;
mem_k_index[7305] = 34262;
mem_k_index[7306] = 34265;
mem_k_index[7307] = 34267;
mem_k_index[7308] = 34270;
mem_k_index[7309] = 34272;
mem_k_index[7310] = 34275;
mem_k_index[7311] = 34277;
mem_k_index[7312] = 34280;
mem_k_index[7313] = 34282;
mem_k_index[7314] = 34285;
mem_k_index[7315] = 34287;
mem_k_index[7316] = 34290;
mem_k_index[7317] = 34292;
mem_k_index[7318] = 34295;
mem_k_index[7319] = 34297;
mem_k_index[7320] = 34300;
mem_k_index[7321] = 34302;
mem_k_index[7322] = 34305;
mem_k_index[7323] = 34307;
mem_k_index[7324] = 34310;
mem_k_index[7325] = 34312;
mem_k_index[7326] = 34315;
mem_k_index[7327] = 34317;
mem_k_index[7328] = 34320;
mem_k_index[7329] = 34322;
mem_k_index[7330] = 34325;
mem_k_index[7331] = 34327;
mem_k_index[7332] = 34330;
mem_k_index[7333] = 34332;
mem_k_index[7334] = 34335;
mem_k_index[7335] = 34337;
mem_k_index[7336] = 34340;
mem_k_index[7337] = 34342;
mem_k_index[7338] = 34345;
mem_k_index[7339] = 34348;
mem_k_index[7340] = 34350;
mem_k_index[7341] = 34353;
mem_k_index[7342] = 34355;
mem_k_index[7343] = 34358;
mem_k_index[7344] = 34360;
mem_k_index[7345] = 34363;
mem_k_index[7346] = 34365;
mem_k_index[7347] = 34368;
mem_k_index[7348] = 34370;
mem_k_index[7349] = 34373;
mem_k_index[7350] = 34375;
mem_k_index[7351] = 34378;
mem_k_index[7352] = 34380;
mem_k_index[7353] = 34383;
mem_k_index[7354] = 34385;
mem_k_index[7355] = 34388;
mem_k_index[7356] = 34390;
mem_k_index[7357] = 34393;
mem_k_index[7358] = 34395;
mem_k_index[7359] = 34398;
mem_k_index[7360] = 34400;
mem_k_index[7361] = 34403;
mem_k_index[7362] = 34405;
mem_k_index[7363] = 34408;
mem_k_index[7364] = 34410;
mem_k_index[7365] = 34413;
mem_k_index[7366] = 34415;
mem_k_index[7367] = 34418;
mem_k_index[7368] = 34420;
mem_k_index[7369] = 34423;
mem_k_index[7370] = 34425;
mem_k_index[7371] = 34428;
mem_k_index[7372] = 34430;
mem_k_index[7373] = 34433;
mem_k_index[7374] = 34435;
mem_k_index[7375] = 34438;
mem_k_index[7376] = 34440;
mem_k_index[7377] = 34443;
mem_k_index[7378] = 34445;
mem_k_index[7379] = 34448;
mem_k_index[7380] = 34450;
mem_k_index[7381] = 34453;
mem_k_index[7382] = 34456;
mem_k_index[7383] = 34458;
mem_k_index[7384] = 34461;
mem_k_index[7385] = 34463;
mem_k_index[7386] = 34466;
mem_k_index[7387] = 34468;
mem_k_index[7388] = 34471;
mem_k_index[7389] = 34473;
mem_k_index[7390] = 34476;
mem_k_index[7391] = 34478;
mem_k_index[7392] = 34481;
mem_k_index[7393] = 34483;
mem_k_index[7394] = 34486;
mem_k_index[7395] = 34488;
mem_k_index[7396] = 34491;
mem_k_index[7397] = 34493;
mem_k_index[7398] = 34496;
mem_k_index[7399] = 34498;
mem_k_index[7400] = 34501;
mem_k_index[7401] = 34503;
mem_k_index[7402] = 34506;
mem_k_index[7403] = 34508;
mem_k_index[7404] = 34511;
mem_k_index[7405] = 34513;
mem_k_index[7406] = 34516;
mem_k_index[7407] = 34518;
mem_k_index[7408] = 34521;
mem_k_index[7409] = 34523;
mem_k_index[7410] = 34526;
mem_k_index[7411] = 34528;
mem_k_index[7412] = 34531;
mem_k_index[7413] = 34533;
mem_k_index[7414] = 34536;
mem_k_index[7415] = 34538;
mem_k_index[7416] = 34541;
mem_k_index[7417] = 34543;
mem_k_index[7418] = 34546;
mem_k_index[7419] = 34548;
mem_k_index[7420] = 34551;
mem_k_index[7421] = 34553;
mem_k_index[7422] = 34556;
mem_k_index[7423] = 34558;
mem_k_index[7424] = 34880;
mem_k_index[7425] = 34882;
mem_k_index[7426] = 34885;
mem_k_index[7427] = 34887;
mem_k_index[7428] = 34890;
mem_k_index[7429] = 34892;
mem_k_index[7430] = 34895;
mem_k_index[7431] = 34897;
mem_k_index[7432] = 34900;
mem_k_index[7433] = 34902;
mem_k_index[7434] = 34905;
mem_k_index[7435] = 34907;
mem_k_index[7436] = 34910;
mem_k_index[7437] = 34912;
mem_k_index[7438] = 34915;
mem_k_index[7439] = 34917;
mem_k_index[7440] = 34920;
mem_k_index[7441] = 34922;
mem_k_index[7442] = 34925;
mem_k_index[7443] = 34927;
mem_k_index[7444] = 34930;
mem_k_index[7445] = 34932;
mem_k_index[7446] = 34935;
mem_k_index[7447] = 34937;
mem_k_index[7448] = 34940;
mem_k_index[7449] = 34942;
mem_k_index[7450] = 34945;
mem_k_index[7451] = 34947;
mem_k_index[7452] = 34950;
mem_k_index[7453] = 34952;
mem_k_index[7454] = 34955;
mem_k_index[7455] = 34957;
mem_k_index[7456] = 34960;
mem_k_index[7457] = 34962;
mem_k_index[7458] = 34965;
mem_k_index[7459] = 34967;
mem_k_index[7460] = 34970;
mem_k_index[7461] = 34972;
mem_k_index[7462] = 34975;
mem_k_index[7463] = 34977;
mem_k_index[7464] = 34980;
mem_k_index[7465] = 34982;
mem_k_index[7466] = 34985;
mem_k_index[7467] = 34988;
mem_k_index[7468] = 34990;
mem_k_index[7469] = 34993;
mem_k_index[7470] = 34995;
mem_k_index[7471] = 34998;
mem_k_index[7472] = 35000;
mem_k_index[7473] = 35003;
mem_k_index[7474] = 35005;
mem_k_index[7475] = 35008;
mem_k_index[7476] = 35010;
mem_k_index[7477] = 35013;
mem_k_index[7478] = 35015;
mem_k_index[7479] = 35018;
mem_k_index[7480] = 35020;
mem_k_index[7481] = 35023;
mem_k_index[7482] = 35025;
mem_k_index[7483] = 35028;
mem_k_index[7484] = 35030;
mem_k_index[7485] = 35033;
mem_k_index[7486] = 35035;
mem_k_index[7487] = 35038;
mem_k_index[7488] = 35040;
mem_k_index[7489] = 35043;
mem_k_index[7490] = 35045;
mem_k_index[7491] = 35048;
mem_k_index[7492] = 35050;
mem_k_index[7493] = 35053;
mem_k_index[7494] = 35055;
mem_k_index[7495] = 35058;
mem_k_index[7496] = 35060;
mem_k_index[7497] = 35063;
mem_k_index[7498] = 35065;
mem_k_index[7499] = 35068;
mem_k_index[7500] = 35070;
mem_k_index[7501] = 35073;
mem_k_index[7502] = 35075;
mem_k_index[7503] = 35078;
mem_k_index[7504] = 35080;
mem_k_index[7505] = 35083;
mem_k_index[7506] = 35085;
mem_k_index[7507] = 35088;
mem_k_index[7508] = 35090;
mem_k_index[7509] = 35093;
mem_k_index[7510] = 35096;
mem_k_index[7511] = 35098;
mem_k_index[7512] = 35101;
mem_k_index[7513] = 35103;
mem_k_index[7514] = 35106;
mem_k_index[7515] = 35108;
mem_k_index[7516] = 35111;
mem_k_index[7517] = 35113;
mem_k_index[7518] = 35116;
mem_k_index[7519] = 35118;
mem_k_index[7520] = 35121;
mem_k_index[7521] = 35123;
mem_k_index[7522] = 35126;
mem_k_index[7523] = 35128;
mem_k_index[7524] = 35131;
mem_k_index[7525] = 35133;
mem_k_index[7526] = 35136;
mem_k_index[7527] = 35138;
mem_k_index[7528] = 35141;
mem_k_index[7529] = 35143;
mem_k_index[7530] = 35146;
mem_k_index[7531] = 35148;
mem_k_index[7532] = 35151;
mem_k_index[7533] = 35153;
mem_k_index[7534] = 35156;
mem_k_index[7535] = 35158;
mem_k_index[7536] = 35161;
mem_k_index[7537] = 35163;
mem_k_index[7538] = 35166;
mem_k_index[7539] = 35168;
mem_k_index[7540] = 35171;
mem_k_index[7541] = 35173;
mem_k_index[7542] = 35176;
mem_k_index[7543] = 35178;
mem_k_index[7544] = 35181;
mem_k_index[7545] = 35183;
mem_k_index[7546] = 35186;
mem_k_index[7547] = 35188;
mem_k_index[7548] = 35191;
mem_k_index[7549] = 35193;
mem_k_index[7550] = 35196;
mem_k_index[7551] = 35198;
mem_k_index[7552] = 35520;
mem_k_index[7553] = 35522;
mem_k_index[7554] = 35525;
mem_k_index[7555] = 35527;
mem_k_index[7556] = 35530;
mem_k_index[7557] = 35532;
mem_k_index[7558] = 35535;
mem_k_index[7559] = 35537;
mem_k_index[7560] = 35540;
mem_k_index[7561] = 35542;
mem_k_index[7562] = 35545;
mem_k_index[7563] = 35547;
mem_k_index[7564] = 35550;
mem_k_index[7565] = 35552;
mem_k_index[7566] = 35555;
mem_k_index[7567] = 35557;
mem_k_index[7568] = 35560;
mem_k_index[7569] = 35562;
mem_k_index[7570] = 35565;
mem_k_index[7571] = 35567;
mem_k_index[7572] = 35570;
mem_k_index[7573] = 35572;
mem_k_index[7574] = 35575;
mem_k_index[7575] = 35577;
mem_k_index[7576] = 35580;
mem_k_index[7577] = 35582;
mem_k_index[7578] = 35585;
mem_k_index[7579] = 35587;
mem_k_index[7580] = 35590;
mem_k_index[7581] = 35592;
mem_k_index[7582] = 35595;
mem_k_index[7583] = 35597;
mem_k_index[7584] = 35600;
mem_k_index[7585] = 35602;
mem_k_index[7586] = 35605;
mem_k_index[7587] = 35607;
mem_k_index[7588] = 35610;
mem_k_index[7589] = 35612;
mem_k_index[7590] = 35615;
mem_k_index[7591] = 35617;
mem_k_index[7592] = 35620;
mem_k_index[7593] = 35622;
mem_k_index[7594] = 35625;
mem_k_index[7595] = 35628;
mem_k_index[7596] = 35630;
mem_k_index[7597] = 35633;
mem_k_index[7598] = 35635;
mem_k_index[7599] = 35638;
mem_k_index[7600] = 35640;
mem_k_index[7601] = 35643;
mem_k_index[7602] = 35645;
mem_k_index[7603] = 35648;
mem_k_index[7604] = 35650;
mem_k_index[7605] = 35653;
mem_k_index[7606] = 35655;
mem_k_index[7607] = 35658;
mem_k_index[7608] = 35660;
mem_k_index[7609] = 35663;
mem_k_index[7610] = 35665;
mem_k_index[7611] = 35668;
mem_k_index[7612] = 35670;
mem_k_index[7613] = 35673;
mem_k_index[7614] = 35675;
mem_k_index[7615] = 35678;
mem_k_index[7616] = 35680;
mem_k_index[7617] = 35683;
mem_k_index[7618] = 35685;
mem_k_index[7619] = 35688;
mem_k_index[7620] = 35690;
mem_k_index[7621] = 35693;
mem_k_index[7622] = 35695;
mem_k_index[7623] = 35698;
mem_k_index[7624] = 35700;
mem_k_index[7625] = 35703;
mem_k_index[7626] = 35705;
mem_k_index[7627] = 35708;
mem_k_index[7628] = 35710;
mem_k_index[7629] = 35713;
mem_k_index[7630] = 35715;
mem_k_index[7631] = 35718;
mem_k_index[7632] = 35720;
mem_k_index[7633] = 35723;
mem_k_index[7634] = 35725;
mem_k_index[7635] = 35728;
mem_k_index[7636] = 35730;
mem_k_index[7637] = 35733;
mem_k_index[7638] = 35736;
mem_k_index[7639] = 35738;
mem_k_index[7640] = 35741;
mem_k_index[7641] = 35743;
mem_k_index[7642] = 35746;
mem_k_index[7643] = 35748;
mem_k_index[7644] = 35751;
mem_k_index[7645] = 35753;
mem_k_index[7646] = 35756;
mem_k_index[7647] = 35758;
mem_k_index[7648] = 35761;
mem_k_index[7649] = 35763;
mem_k_index[7650] = 35766;
mem_k_index[7651] = 35768;
mem_k_index[7652] = 35771;
mem_k_index[7653] = 35773;
mem_k_index[7654] = 35776;
mem_k_index[7655] = 35778;
mem_k_index[7656] = 35781;
mem_k_index[7657] = 35783;
mem_k_index[7658] = 35786;
mem_k_index[7659] = 35788;
mem_k_index[7660] = 35791;
mem_k_index[7661] = 35793;
mem_k_index[7662] = 35796;
mem_k_index[7663] = 35798;
mem_k_index[7664] = 35801;
mem_k_index[7665] = 35803;
mem_k_index[7666] = 35806;
mem_k_index[7667] = 35808;
mem_k_index[7668] = 35811;
mem_k_index[7669] = 35813;
mem_k_index[7670] = 35816;
mem_k_index[7671] = 35818;
mem_k_index[7672] = 35821;
mem_k_index[7673] = 35823;
mem_k_index[7674] = 35826;
mem_k_index[7675] = 35828;
mem_k_index[7676] = 35831;
mem_k_index[7677] = 35833;
mem_k_index[7678] = 35836;
mem_k_index[7679] = 35838;
mem_k_index[7680] = 35840;
mem_k_index[7681] = 35842;
mem_k_index[7682] = 35845;
mem_k_index[7683] = 35847;
mem_k_index[7684] = 35850;
mem_k_index[7685] = 35852;
mem_k_index[7686] = 35855;
mem_k_index[7687] = 35857;
mem_k_index[7688] = 35860;
mem_k_index[7689] = 35862;
mem_k_index[7690] = 35865;
mem_k_index[7691] = 35867;
mem_k_index[7692] = 35870;
mem_k_index[7693] = 35872;
mem_k_index[7694] = 35875;
mem_k_index[7695] = 35877;
mem_k_index[7696] = 35880;
mem_k_index[7697] = 35882;
mem_k_index[7698] = 35885;
mem_k_index[7699] = 35887;
mem_k_index[7700] = 35890;
mem_k_index[7701] = 35892;
mem_k_index[7702] = 35895;
mem_k_index[7703] = 35897;
mem_k_index[7704] = 35900;
mem_k_index[7705] = 35902;
mem_k_index[7706] = 35905;
mem_k_index[7707] = 35907;
mem_k_index[7708] = 35910;
mem_k_index[7709] = 35912;
mem_k_index[7710] = 35915;
mem_k_index[7711] = 35917;
mem_k_index[7712] = 35920;
mem_k_index[7713] = 35922;
mem_k_index[7714] = 35925;
mem_k_index[7715] = 35927;
mem_k_index[7716] = 35930;
mem_k_index[7717] = 35932;
mem_k_index[7718] = 35935;
mem_k_index[7719] = 35937;
mem_k_index[7720] = 35940;
mem_k_index[7721] = 35942;
mem_k_index[7722] = 35945;
mem_k_index[7723] = 35948;
mem_k_index[7724] = 35950;
mem_k_index[7725] = 35953;
mem_k_index[7726] = 35955;
mem_k_index[7727] = 35958;
mem_k_index[7728] = 35960;
mem_k_index[7729] = 35963;
mem_k_index[7730] = 35965;
mem_k_index[7731] = 35968;
mem_k_index[7732] = 35970;
mem_k_index[7733] = 35973;
mem_k_index[7734] = 35975;
mem_k_index[7735] = 35978;
mem_k_index[7736] = 35980;
mem_k_index[7737] = 35983;
mem_k_index[7738] = 35985;
mem_k_index[7739] = 35988;
mem_k_index[7740] = 35990;
mem_k_index[7741] = 35993;
mem_k_index[7742] = 35995;
mem_k_index[7743] = 35998;
mem_k_index[7744] = 36000;
mem_k_index[7745] = 36003;
mem_k_index[7746] = 36005;
mem_k_index[7747] = 36008;
mem_k_index[7748] = 36010;
mem_k_index[7749] = 36013;
mem_k_index[7750] = 36015;
mem_k_index[7751] = 36018;
mem_k_index[7752] = 36020;
mem_k_index[7753] = 36023;
mem_k_index[7754] = 36025;
mem_k_index[7755] = 36028;
mem_k_index[7756] = 36030;
mem_k_index[7757] = 36033;
mem_k_index[7758] = 36035;
mem_k_index[7759] = 36038;
mem_k_index[7760] = 36040;
mem_k_index[7761] = 36043;
mem_k_index[7762] = 36045;
mem_k_index[7763] = 36048;
mem_k_index[7764] = 36050;
mem_k_index[7765] = 36053;
mem_k_index[7766] = 36056;
mem_k_index[7767] = 36058;
mem_k_index[7768] = 36061;
mem_k_index[7769] = 36063;
mem_k_index[7770] = 36066;
mem_k_index[7771] = 36068;
mem_k_index[7772] = 36071;
mem_k_index[7773] = 36073;
mem_k_index[7774] = 36076;
mem_k_index[7775] = 36078;
mem_k_index[7776] = 36081;
mem_k_index[7777] = 36083;
mem_k_index[7778] = 36086;
mem_k_index[7779] = 36088;
mem_k_index[7780] = 36091;
mem_k_index[7781] = 36093;
mem_k_index[7782] = 36096;
mem_k_index[7783] = 36098;
mem_k_index[7784] = 36101;
mem_k_index[7785] = 36103;
mem_k_index[7786] = 36106;
mem_k_index[7787] = 36108;
mem_k_index[7788] = 36111;
mem_k_index[7789] = 36113;
mem_k_index[7790] = 36116;
mem_k_index[7791] = 36118;
mem_k_index[7792] = 36121;
mem_k_index[7793] = 36123;
mem_k_index[7794] = 36126;
mem_k_index[7795] = 36128;
mem_k_index[7796] = 36131;
mem_k_index[7797] = 36133;
mem_k_index[7798] = 36136;
mem_k_index[7799] = 36138;
mem_k_index[7800] = 36141;
mem_k_index[7801] = 36143;
mem_k_index[7802] = 36146;
mem_k_index[7803] = 36148;
mem_k_index[7804] = 36151;
mem_k_index[7805] = 36153;
mem_k_index[7806] = 36156;
mem_k_index[7807] = 36158;
mem_k_index[7808] = 36480;
mem_k_index[7809] = 36482;
mem_k_index[7810] = 36485;
mem_k_index[7811] = 36487;
mem_k_index[7812] = 36490;
mem_k_index[7813] = 36492;
mem_k_index[7814] = 36495;
mem_k_index[7815] = 36497;
mem_k_index[7816] = 36500;
mem_k_index[7817] = 36502;
mem_k_index[7818] = 36505;
mem_k_index[7819] = 36507;
mem_k_index[7820] = 36510;
mem_k_index[7821] = 36512;
mem_k_index[7822] = 36515;
mem_k_index[7823] = 36517;
mem_k_index[7824] = 36520;
mem_k_index[7825] = 36522;
mem_k_index[7826] = 36525;
mem_k_index[7827] = 36527;
mem_k_index[7828] = 36530;
mem_k_index[7829] = 36532;
mem_k_index[7830] = 36535;
mem_k_index[7831] = 36537;
mem_k_index[7832] = 36540;
mem_k_index[7833] = 36542;
mem_k_index[7834] = 36545;
mem_k_index[7835] = 36547;
mem_k_index[7836] = 36550;
mem_k_index[7837] = 36552;
mem_k_index[7838] = 36555;
mem_k_index[7839] = 36557;
mem_k_index[7840] = 36560;
mem_k_index[7841] = 36562;
mem_k_index[7842] = 36565;
mem_k_index[7843] = 36567;
mem_k_index[7844] = 36570;
mem_k_index[7845] = 36572;
mem_k_index[7846] = 36575;
mem_k_index[7847] = 36577;
mem_k_index[7848] = 36580;
mem_k_index[7849] = 36582;
mem_k_index[7850] = 36585;
mem_k_index[7851] = 36588;
mem_k_index[7852] = 36590;
mem_k_index[7853] = 36593;
mem_k_index[7854] = 36595;
mem_k_index[7855] = 36598;
mem_k_index[7856] = 36600;
mem_k_index[7857] = 36603;
mem_k_index[7858] = 36605;
mem_k_index[7859] = 36608;
mem_k_index[7860] = 36610;
mem_k_index[7861] = 36613;
mem_k_index[7862] = 36615;
mem_k_index[7863] = 36618;
mem_k_index[7864] = 36620;
mem_k_index[7865] = 36623;
mem_k_index[7866] = 36625;
mem_k_index[7867] = 36628;
mem_k_index[7868] = 36630;
mem_k_index[7869] = 36633;
mem_k_index[7870] = 36635;
mem_k_index[7871] = 36638;
mem_k_index[7872] = 36640;
mem_k_index[7873] = 36643;
mem_k_index[7874] = 36645;
mem_k_index[7875] = 36648;
mem_k_index[7876] = 36650;
mem_k_index[7877] = 36653;
mem_k_index[7878] = 36655;
mem_k_index[7879] = 36658;
mem_k_index[7880] = 36660;
mem_k_index[7881] = 36663;
mem_k_index[7882] = 36665;
mem_k_index[7883] = 36668;
mem_k_index[7884] = 36670;
mem_k_index[7885] = 36673;
mem_k_index[7886] = 36675;
mem_k_index[7887] = 36678;
mem_k_index[7888] = 36680;
mem_k_index[7889] = 36683;
mem_k_index[7890] = 36685;
mem_k_index[7891] = 36688;
mem_k_index[7892] = 36690;
mem_k_index[7893] = 36693;
mem_k_index[7894] = 36696;
mem_k_index[7895] = 36698;
mem_k_index[7896] = 36701;
mem_k_index[7897] = 36703;
mem_k_index[7898] = 36706;
mem_k_index[7899] = 36708;
mem_k_index[7900] = 36711;
mem_k_index[7901] = 36713;
mem_k_index[7902] = 36716;
mem_k_index[7903] = 36718;
mem_k_index[7904] = 36721;
mem_k_index[7905] = 36723;
mem_k_index[7906] = 36726;
mem_k_index[7907] = 36728;
mem_k_index[7908] = 36731;
mem_k_index[7909] = 36733;
mem_k_index[7910] = 36736;
mem_k_index[7911] = 36738;
mem_k_index[7912] = 36741;
mem_k_index[7913] = 36743;
mem_k_index[7914] = 36746;
mem_k_index[7915] = 36748;
mem_k_index[7916] = 36751;
mem_k_index[7917] = 36753;
mem_k_index[7918] = 36756;
mem_k_index[7919] = 36758;
mem_k_index[7920] = 36761;
mem_k_index[7921] = 36763;
mem_k_index[7922] = 36766;
mem_k_index[7923] = 36768;
mem_k_index[7924] = 36771;
mem_k_index[7925] = 36773;
mem_k_index[7926] = 36776;
mem_k_index[7927] = 36778;
mem_k_index[7928] = 36781;
mem_k_index[7929] = 36783;
mem_k_index[7930] = 36786;
mem_k_index[7931] = 36788;
mem_k_index[7932] = 36791;
mem_k_index[7933] = 36793;
mem_k_index[7934] = 36796;
mem_k_index[7935] = 36798;
mem_k_index[7936] = 37120;
mem_k_index[7937] = 37122;
mem_k_index[7938] = 37125;
mem_k_index[7939] = 37127;
mem_k_index[7940] = 37130;
mem_k_index[7941] = 37132;
mem_k_index[7942] = 37135;
mem_k_index[7943] = 37137;
mem_k_index[7944] = 37140;
mem_k_index[7945] = 37142;
mem_k_index[7946] = 37145;
mem_k_index[7947] = 37147;
mem_k_index[7948] = 37150;
mem_k_index[7949] = 37152;
mem_k_index[7950] = 37155;
mem_k_index[7951] = 37157;
mem_k_index[7952] = 37160;
mem_k_index[7953] = 37162;
mem_k_index[7954] = 37165;
mem_k_index[7955] = 37167;
mem_k_index[7956] = 37170;
mem_k_index[7957] = 37172;
mem_k_index[7958] = 37175;
mem_k_index[7959] = 37177;
mem_k_index[7960] = 37180;
mem_k_index[7961] = 37182;
mem_k_index[7962] = 37185;
mem_k_index[7963] = 37187;
mem_k_index[7964] = 37190;
mem_k_index[7965] = 37192;
mem_k_index[7966] = 37195;
mem_k_index[7967] = 37197;
mem_k_index[7968] = 37200;
mem_k_index[7969] = 37202;
mem_k_index[7970] = 37205;
mem_k_index[7971] = 37207;
mem_k_index[7972] = 37210;
mem_k_index[7973] = 37212;
mem_k_index[7974] = 37215;
mem_k_index[7975] = 37217;
mem_k_index[7976] = 37220;
mem_k_index[7977] = 37222;
mem_k_index[7978] = 37225;
mem_k_index[7979] = 37228;
mem_k_index[7980] = 37230;
mem_k_index[7981] = 37233;
mem_k_index[7982] = 37235;
mem_k_index[7983] = 37238;
mem_k_index[7984] = 37240;
mem_k_index[7985] = 37243;
mem_k_index[7986] = 37245;
mem_k_index[7987] = 37248;
mem_k_index[7988] = 37250;
mem_k_index[7989] = 37253;
mem_k_index[7990] = 37255;
mem_k_index[7991] = 37258;
mem_k_index[7992] = 37260;
mem_k_index[7993] = 37263;
mem_k_index[7994] = 37265;
mem_k_index[7995] = 37268;
mem_k_index[7996] = 37270;
mem_k_index[7997] = 37273;
mem_k_index[7998] = 37275;
mem_k_index[7999] = 37278;
mem_k_index[8000] = 37280;
mem_k_index[8001] = 37283;
mem_k_index[8002] = 37285;
mem_k_index[8003] = 37288;
mem_k_index[8004] = 37290;
mem_k_index[8005] = 37293;
mem_k_index[8006] = 37295;
mem_k_index[8007] = 37298;
mem_k_index[8008] = 37300;
mem_k_index[8009] = 37303;
mem_k_index[8010] = 37305;
mem_k_index[8011] = 37308;
mem_k_index[8012] = 37310;
mem_k_index[8013] = 37313;
mem_k_index[8014] = 37315;
mem_k_index[8015] = 37318;
mem_k_index[8016] = 37320;
mem_k_index[8017] = 37323;
mem_k_index[8018] = 37325;
mem_k_index[8019] = 37328;
mem_k_index[8020] = 37330;
mem_k_index[8021] = 37333;
mem_k_index[8022] = 37336;
mem_k_index[8023] = 37338;
mem_k_index[8024] = 37341;
mem_k_index[8025] = 37343;
mem_k_index[8026] = 37346;
mem_k_index[8027] = 37348;
mem_k_index[8028] = 37351;
mem_k_index[8029] = 37353;
mem_k_index[8030] = 37356;
mem_k_index[8031] = 37358;
mem_k_index[8032] = 37361;
mem_k_index[8033] = 37363;
mem_k_index[8034] = 37366;
mem_k_index[8035] = 37368;
mem_k_index[8036] = 37371;
mem_k_index[8037] = 37373;
mem_k_index[8038] = 37376;
mem_k_index[8039] = 37378;
mem_k_index[8040] = 37381;
mem_k_index[8041] = 37383;
mem_k_index[8042] = 37386;
mem_k_index[8043] = 37388;
mem_k_index[8044] = 37391;
mem_k_index[8045] = 37393;
mem_k_index[8046] = 37396;
mem_k_index[8047] = 37398;
mem_k_index[8048] = 37401;
mem_k_index[8049] = 37403;
mem_k_index[8050] = 37406;
mem_k_index[8051] = 37408;
mem_k_index[8052] = 37411;
mem_k_index[8053] = 37413;
mem_k_index[8054] = 37416;
mem_k_index[8055] = 37418;
mem_k_index[8056] = 37421;
mem_k_index[8057] = 37423;
mem_k_index[8058] = 37426;
mem_k_index[8059] = 37428;
mem_k_index[8060] = 37431;
mem_k_index[8061] = 37433;
mem_k_index[8062] = 37436;
mem_k_index[8063] = 37438;
mem_k_index[8064] = 37760;
mem_k_index[8065] = 37762;
mem_k_index[8066] = 37765;
mem_k_index[8067] = 37767;
mem_k_index[8068] = 37770;
mem_k_index[8069] = 37772;
mem_k_index[8070] = 37775;
mem_k_index[8071] = 37777;
mem_k_index[8072] = 37780;
mem_k_index[8073] = 37782;
mem_k_index[8074] = 37785;
mem_k_index[8075] = 37787;
mem_k_index[8076] = 37790;
mem_k_index[8077] = 37792;
mem_k_index[8078] = 37795;
mem_k_index[8079] = 37797;
mem_k_index[8080] = 37800;
mem_k_index[8081] = 37802;
mem_k_index[8082] = 37805;
mem_k_index[8083] = 37807;
mem_k_index[8084] = 37810;
mem_k_index[8085] = 37812;
mem_k_index[8086] = 37815;
mem_k_index[8087] = 37817;
mem_k_index[8088] = 37820;
mem_k_index[8089] = 37822;
mem_k_index[8090] = 37825;
mem_k_index[8091] = 37827;
mem_k_index[8092] = 37830;
mem_k_index[8093] = 37832;
mem_k_index[8094] = 37835;
mem_k_index[8095] = 37837;
mem_k_index[8096] = 37840;
mem_k_index[8097] = 37842;
mem_k_index[8098] = 37845;
mem_k_index[8099] = 37847;
mem_k_index[8100] = 37850;
mem_k_index[8101] = 37852;
mem_k_index[8102] = 37855;
mem_k_index[8103] = 37857;
mem_k_index[8104] = 37860;
mem_k_index[8105] = 37862;
mem_k_index[8106] = 37865;
mem_k_index[8107] = 37868;
mem_k_index[8108] = 37870;
mem_k_index[8109] = 37873;
mem_k_index[8110] = 37875;
mem_k_index[8111] = 37878;
mem_k_index[8112] = 37880;
mem_k_index[8113] = 37883;
mem_k_index[8114] = 37885;
mem_k_index[8115] = 37888;
mem_k_index[8116] = 37890;
mem_k_index[8117] = 37893;
mem_k_index[8118] = 37895;
mem_k_index[8119] = 37898;
mem_k_index[8120] = 37900;
mem_k_index[8121] = 37903;
mem_k_index[8122] = 37905;
mem_k_index[8123] = 37908;
mem_k_index[8124] = 37910;
mem_k_index[8125] = 37913;
mem_k_index[8126] = 37915;
mem_k_index[8127] = 37918;
mem_k_index[8128] = 37920;
mem_k_index[8129] = 37923;
mem_k_index[8130] = 37925;
mem_k_index[8131] = 37928;
mem_k_index[8132] = 37930;
mem_k_index[8133] = 37933;
mem_k_index[8134] = 37935;
mem_k_index[8135] = 37938;
mem_k_index[8136] = 37940;
mem_k_index[8137] = 37943;
mem_k_index[8138] = 37945;
mem_k_index[8139] = 37948;
mem_k_index[8140] = 37950;
mem_k_index[8141] = 37953;
mem_k_index[8142] = 37955;
mem_k_index[8143] = 37958;
mem_k_index[8144] = 37960;
mem_k_index[8145] = 37963;
mem_k_index[8146] = 37965;
mem_k_index[8147] = 37968;
mem_k_index[8148] = 37970;
mem_k_index[8149] = 37973;
mem_k_index[8150] = 37976;
mem_k_index[8151] = 37978;
mem_k_index[8152] = 37981;
mem_k_index[8153] = 37983;
mem_k_index[8154] = 37986;
mem_k_index[8155] = 37988;
mem_k_index[8156] = 37991;
mem_k_index[8157] = 37993;
mem_k_index[8158] = 37996;
mem_k_index[8159] = 37998;
mem_k_index[8160] = 38001;
mem_k_index[8161] = 38003;
mem_k_index[8162] = 38006;
mem_k_index[8163] = 38008;
mem_k_index[8164] = 38011;
mem_k_index[8165] = 38013;
mem_k_index[8166] = 38016;
mem_k_index[8167] = 38018;
mem_k_index[8168] = 38021;
mem_k_index[8169] = 38023;
mem_k_index[8170] = 38026;
mem_k_index[8171] = 38028;
mem_k_index[8172] = 38031;
mem_k_index[8173] = 38033;
mem_k_index[8174] = 38036;
mem_k_index[8175] = 38038;
mem_k_index[8176] = 38041;
mem_k_index[8177] = 38043;
mem_k_index[8178] = 38046;
mem_k_index[8179] = 38048;
mem_k_index[8180] = 38051;
mem_k_index[8181] = 38053;
mem_k_index[8182] = 38056;
mem_k_index[8183] = 38058;
mem_k_index[8184] = 38061;
mem_k_index[8185] = 38063;
mem_k_index[8186] = 38066;
mem_k_index[8187] = 38068;
mem_k_index[8188] = 38071;
mem_k_index[8189] = 38073;
mem_k_index[8190] = 38076;
mem_k_index[8191] = 38078;
mem_k_index[8192] = 38400;
mem_k_index[8193] = 38402;
mem_k_index[8194] = 38405;
mem_k_index[8195] = 38407;
mem_k_index[8196] = 38410;
mem_k_index[8197] = 38412;
mem_k_index[8198] = 38415;
mem_k_index[8199] = 38417;
mem_k_index[8200] = 38420;
mem_k_index[8201] = 38422;
mem_k_index[8202] = 38425;
mem_k_index[8203] = 38427;
mem_k_index[8204] = 38430;
mem_k_index[8205] = 38432;
mem_k_index[8206] = 38435;
mem_k_index[8207] = 38437;
mem_k_index[8208] = 38440;
mem_k_index[8209] = 38442;
mem_k_index[8210] = 38445;
mem_k_index[8211] = 38447;
mem_k_index[8212] = 38450;
mem_k_index[8213] = 38452;
mem_k_index[8214] = 38455;
mem_k_index[8215] = 38457;
mem_k_index[8216] = 38460;
mem_k_index[8217] = 38462;
mem_k_index[8218] = 38465;
mem_k_index[8219] = 38467;
mem_k_index[8220] = 38470;
mem_k_index[8221] = 38472;
mem_k_index[8222] = 38475;
mem_k_index[8223] = 38477;
mem_k_index[8224] = 38480;
mem_k_index[8225] = 38482;
mem_k_index[8226] = 38485;
mem_k_index[8227] = 38487;
mem_k_index[8228] = 38490;
mem_k_index[8229] = 38492;
mem_k_index[8230] = 38495;
mem_k_index[8231] = 38497;
mem_k_index[8232] = 38500;
mem_k_index[8233] = 38502;
mem_k_index[8234] = 38505;
mem_k_index[8235] = 38508;
mem_k_index[8236] = 38510;
mem_k_index[8237] = 38513;
mem_k_index[8238] = 38515;
mem_k_index[8239] = 38518;
mem_k_index[8240] = 38520;
mem_k_index[8241] = 38523;
mem_k_index[8242] = 38525;
mem_k_index[8243] = 38528;
mem_k_index[8244] = 38530;
mem_k_index[8245] = 38533;
mem_k_index[8246] = 38535;
mem_k_index[8247] = 38538;
mem_k_index[8248] = 38540;
mem_k_index[8249] = 38543;
mem_k_index[8250] = 38545;
mem_k_index[8251] = 38548;
mem_k_index[8252] = 38550;
mem_k_index[8253] = 38553;
mem_k_index[8254] = 38555;
mem_k_index[8255] = 38558;
mem_k_index[8256] = 38560;
mem_k_index[8257] = 38563;
mem_k_index[8258] = 38565;
mem_k_index[8259] = 38568;
mem_k_index[8260] = 38570;
mem_k_index[8261] = 38573;
mem_k_index[8262] = 38575;
mem_k_index[8263] = 38578;
mem_k_index[8264] = 38580;
mem_k_index[8265] = 38583;
mem_k_index[8266] = 38585;
mem_k_index[8267] = 38588;
mem_k_index[8268] = 38590;
mem_k_index[8269] = 38593;
mem_k_index[8270] = 38595;
mem_k_index[8271] = 38598;
mem_k_index[8272] = 38600;
mem_k_index[8273] = 38603;
mem_k_index[8274] = 38605;
mem_k_index[8275] = 38608;
mem_k_index[8276] = 38610;
mem_k_index[8277] = 38613;
mem_k_index[8278] = 38616;
mem_k_index[8279] = 38618;
mem_k_index[8280] = 38621;
mem_k_index[8281] = 38623;
mem_k_index[8282] = 38626;
mem_k_index[8283] = 38628;
mem_k_index[8284] = 38631;
mem_k_index[8285] = 38633;
mem_k_index[8286] = 38636;
mem_k_index[8287] = 38638;
mem_k_index[8288] = 38641;
mem_k_index[8289] = 38643;
mem_k_index[8290] = 38646;
mem_k_index[8291] = 38648;
mem_k_index[8292] = 38651;
mem_k_index[8293] = 38653;
mem_k_index[8294] = 38656;
mem_k_index[8295] = 38658;
mem_k_index[8296] = 38661;
mem_k_index[8297] = 38663;
mem_k_index[8298] = 38666;
mem_k_index[8299] = 38668;
mem_k_index[8300] = 38671;
mem_k_index[8301] = 38673;
mem_k_index[8302] = 38676;
mem_k_index[8303] = 38678;
mem_k_index[8304] = 38681;
mem_k_index[8305] = 38683;
mem_k_index[8306] = 38686;
mem_k_index[8307] = 38688;
mem_k_index[8308] = 38691;
mem_k_index[8309] = 38693;
mem_k_index[8310] = 38696;
mem_k_index[8311] = 38698;
mem_k_index[8312] = 38701;
mem_k_index[8313] = 38703;
mem_k_index[8314] = 38706;
mem_k_index[8315] = 38708;
mem_k_index[8316] = 38711;
mem_k_index[8317] = 38713;
mem_k_index[8318] = 38716;
mem_k_index[8319] = 38718;
mem_k_index[8320] = 39040;
mem_k_index[8321] = 39042;
mem_k_index[8322] = 39045;
mem_k_index[8323] = 39047;
mem_k_index[8324] = 39050;
mem_k_index[8325] = 39052;
mem_k_index[8326] = 39055;
mem_k_index[8327] = 39057;
mem_k_index[8328] = 39060;
mem_k_index[8329] = 39062;
mem_k_index[8330] = 39065;
mem_k_index[8331] = 39067;
mem_k_index[8332] = 39070;
mem_k_index[8333] = 39072;
mem_k_index[8334] = 39075;
mem_k_index[8335] = 39077;
mem_k_index[8336] = 39080;
mem_k_index[8337] = 39082;
mem_k_index[8338] = 39085;
mem_k_index[8339] = 39087;
mem_k_index[8340] = 39090;
mem_k_index[8341] = 39092;
mem_k_index[8342] = 39095;
mem_k_index[8343] = 39097;
mem_k_index[8344] = 39100;
mem_k_index[8345] = 39102;
mem_k_index[8346] = 39105;
mem_k_index[8347] = 39107;
mem_k_index[8348] = 39110;
mem_k_index[8349] = 39112;
mem_k_index[8350] = 39115;
mem_k_index[8351] = 39117;
mem_k_index[8352] = 39120;
mem_k_index[8353] = 39122;
mem_k_index[8354] = 39125;
mem_k_index[8355] = 39127;
mem_k_index[8356] = 39130;
mem_k_index[8357] = 39132;
mem_k_index[8358] = 39135;
mem_k_index[8359] = 39137;
mem_k_index[8360] = 39140;
mem_k_index[8361] = 39142;
mem_k_index[8362] = 39145;
mem_k_index[8363] = 39148;
mem_k_index[8364] = 39150;
mem_k_index[8365] = 39153;
mem_k_index[8366] = 39155;
mem_k_index[8367] = 39158;
mem_k_index[8368] = 39160;
mem_k_index[8369] = 39163;
mem_k_index[8370] = 39165;
mem_k_index[8371] = 39168;
mem_k_index[8372] = 39170;
mem_k_index[8373] = 39173;
mem_k_index[8374] = 39175;
mem_k_index[8375] = 39178;
mem_k_index[8376] = 39180;
mem_k_index[8377] = 39183;
mem_k_index[8378] = 39185;
mem_k_index[8379] = 39188;
mem_k_index[8380] = 39190;
mem_k_index[8381] = 39193;
mem_k_index[8382] = 39195;
mem_k_index[8383] = 39198;
mem_k_index[8384] = 39200;
mem_k_index[8385] = 39203;
mem_k_index[8386] = 39205;
mem_k_index[8387] = 39208;
mem_k_index[8388] = 39210;
mem_k_index[8389] = 39213;
mem_k_index[8390] = 39215;
mem_k_index[8391] = 39218;
mem_k_index[8392] = 39220;
mem_k_index[8393] = 39223;
mem_k_index[8394] = 39225;
mem_k_index[8395] = 39228;
mem_k_index[8396] = 39230;
mem_k_index[8397] = 39233;
mem_k_index[8398] = 39235;
mem_k_index[8399] = 39238;
mem_k_index[8400] = 39240;
mem_k_index[8401] = 39243;
mem_k_index[8402] = 39245;
mem_k_index[8403] = 39248;
mem_k_index[8404] = 39250;
mem_k_index[8405] = 39253;
mem_k_index[8406] = 39256;
mem_k_index[8407] = 39258;
mem_k_index[8408] = 39261;
mem_k_index[8409] = 39263;
mem_k_index[8410] = 39266;
mem_k_index[8411] = 39268;
mem_k_index[8412] = 39271;
mem_k_index[8413] = 39273;
mem_k_index[8414] = 39276;
mem_k_index[8415] = 39278;
mem_k_index[8416] = 39281;
mem_k_index[8417] = 39283;
mem_k_index[8418] = 39286;
mem_k_index[8419] = 39288;
mem_k_index[8420] = 39291;
mem_k_index[8421] = 39293;
mem_k_index[8422] = 39296;
mem_k_index[8423] = 39298;
mem_k_index[8424] = 39301;
mem_k_index[8425] = 39303;
mem_k_index[8426] = 39306;
mem_k_index[8427] = 39308;
mem_k_index[8428] = 39311;
mem_k_index[8429] = 39313;
mem_k_index[8430] = 39316;
mem_k_index[8431] = 39318;
mem_k_index[8432] = 39321;
mem_k_index[8433] = 39323;
mem_k_index[8434] = 39326;
mem_k_index[8435] = 39328;
mem_k_index[8436] = 39331;
mem_k_index[8437] = 39333;
mem_k_index[8438] = 39336;
mem_k_index[8439] = 39338;
mem_k_index[8440] = 39341;
mem_k_index[8441] = 39343;
mem_k_index[8442] = 39346;
mem_k_index[8443] = 39348;
mem_k_index[8444] = 39351;
mem_k_index[8445] = 39353;
mem_k_index[8446] = 39356;
mem_k_index[8447] = 39358;
mem_k_index[8448] = 39680;
mem_k_index[8449] = 39682;
mem_k_index[8450] = 39685;
mem_k_index[8451] = 39687;
mem_k_index[8452] = 39690;
mem_k_index[8453] = 39692;
mem_k_index[8454] = 39695;
mem_k_index[8455] = 39697;
mem_k_index[8456] = 39700;
mem_k_index[8457] = 39702;
mem_k_index[8458] = 39705;
mem_k_index[8459] = 39707;
mem_k_index[8460] = 39710;
mem_k_index[8461] = 39712;
mem_k_index[8462] = 39715;
mem_k_index[8463] = 39717;
mem_k_index[8464] = 39720;
mem_k_index[8465] = 39722;
mem_k_index[8466] = 39725;
mem_k_index[8467] = 39727;
mem_k_index[8468] = 39730;
mem_k_index[8469] = 39732;
mem_k_index[8470] = 39735;
mem_k_index[8471] = 39737;
mem_k_index[8472] = 39740;
mem_k_index[8473] = 39742;
mem_k_index[8474] = 39745;
mem_k_index[8475] = 39747;
mem_k_index[8476] = 39750;
mem_k_index[8477] = 39752;
mem_k_index[8478] = 39755;
mem_k_index[8479] = 39757;
mem_k_index[8480] = 39760;
mem_k_index[8481] = 39762;
mem_k_index[8482] = 39765;
mem_k_index[8483] = 39767;
mem_k_index[8484] = 39770;
mem_k_index[8485] = 39772;
mem_k_index[8486] = 39775;
mem_k_index[8487] = 39777;
mem_k_index[8488] = 39780;
mem_k_index[8489] = 39782;
mem_k_index[8490] = 39785;
mem_k_index[8491] = 39788;
mem_k_index[8492] = 39790;
mem_k_index[8493] = 39793;
mem_k_index[8494] = 39795;
mem_k_index[8495] = 39798;
mem_k_index[8496] = 39800;
mem_k_index[8497] = 39803;
mem_k_index[8498] = 39805;
mem_k_index[8499] = 39808;
mem_k_index[8500] = 39810;
mem_k_index[8501] = 39813;
mem_k_index[8502] = 39815;
mem_k_index[8503] = 39818;
mem_k_index[8504] = 39820;
mem_k_index[8505] = 39823;
mem_k_index[8506] = 39825;
mem_k_index[8507] = 39828;
mem_k_index[8508] = 39830;
mem_k_index[8509] = 39833;
mem_k_index[8510] = 39835;
mem_k_index[8511] = 39838;
mem_k_index[8512] = 39840;
mem_k_index[8513] = 39843;
mem_k_index[8514] = 39845;
mem_k_index[8515] = 39848;
mem_k_index[8516] = 39850;
mem_k_index[8517] = 39853;
mem_k_index[8518] = 39855;
mem_k_index[8519] = 39858;
mem_k_index[8520] = 39860;
mem_k_index[8521] = 39863;
mem_k_index[8522] = 39865;
mem_k_index[8523] = 39868;
mem_k_index[8524] = 39870;
mem_k_index[8525] = 39873;
mem_k_index[8526] = 39875;
mem_k_index[8527] = 39878;
mem_k_index[8528] = 39880;
mem_k_index[8529] = 39883;
mem_k_index[8530] = 39885;
mem_k_index[8531] = 39888;
mem_k_index[8532] = 39890;
mem_k_index[8533] = 39893;
mem_k_index[8534] = 39896;
mem_k_index[8535] = 39898;
mem_k_index[8536] = 39901;
mem_k_index[8537] = 39903;
mem_k_index[8538] = 39906;
mem_k_index[8539] = 39908;
mem_k_index[8540] = 39911;
mem_k_index[8541] = 39913;
mem_k_index[8542] = 39916;
mem_k_index[8543] = 39918;
mem_k_index[8544] = 39921;
mem_k_index[8545] = 39923;
mem_k_index[8546] = 39926;
mem_k_index[8547] = 39928;
mem_k_index[8548] = 39931;
mem_k_index[8549] = 39933;
mem_k_index[8550] = 39936;
mem_k_index[8551] = 39938;
mem_k_index[8552] = 39941;
mem_k_index[8553] = 39943;
mem_k_index[8554] = 39946;
mem_k_index[8555] = 39948;
mem_k_index[8556] = 39951;
mem_k_index[8557] = 39953;
mem_k_index[8558] = 39956;
mem_k_index[8559] = 39958;
mem_k_index[8560] = 39961;
mem_k_index[8561] = 39963;
mem_k_index[8562] = 39966;
mem_k_index[8563] = 39968;
mem_k_index[8564] = 39971;
mem_k_index[8565] = 39973;
mem_k_index[8566] = 39976;
mem_k_index[8567] = 39978;
mem_k_index[8568] = 39981;
mem_k_index[8569] = 39983;
mem_k_index[8570] = 39986;
mem_k_index[8571] = 39988;
mem_k_index[8572] = 39991;
mem_k_index[8573] = 39993;
mem_k_index[8574] = 39996;
mem_k_index[8575] = 39998;
mem_k_index[8576] = 40320;
mem_k_index[8577] = 40322;
mem_k_index[8578] = 40325;
mem_k_index[8579] = 40327;
mem_k_index[8580] = 40330;
mem_k_index[8581] = 40332;
mem_k_index[8582] = 40335;
mem_k_index[8583] = 40337;
mem_k_index[8584] = 40340;
mem_k_index[8585] = 40342;
mem_k_index[8586] = 40345;
mem_k_index[8587] = 40347;
mem_k_index[8588] = 40350;
mem_k_index[8589] = 40352;
mem_k_index[8590] = 40355;
mem_k_index[8591] = 40357;
mem_k_index[8592] = 40360;
mem_k_index[8593] = 40362;
mem_k_index[8594] = 40365;
mem_k_index[8595] = 40367;
mem_k_index[8596] = 40370;
mem_k_index[8597] = 40372;
mem_k_index[8598] = 40375;
mem_k_index[8599] = 40377;
mem_k_index[8600] = 40380;
mem_k_index[8601] = 40382;
mem_k_index[8602] = 40385;
mem_k_index[8603] = 40387;
mem_k_index[8604] = 40390;
mem_k_index[8605] = 40392;
mem_k_index[8606] = 40395;
mem_k_index[8607] = 40397;
mem_k_index[8608] = 40400;
mem_k_index[8609] = 40402;
mem_k_index[8610] = 40405;
mem_k_index[8611] = 40407;
mem_k_index[8612] = 40410;
mem_k_index[8613] = 40412;
mem_k_index[8614] = 40415;
mem_k_index[8615] = 40417;
mem_k_index[8616] = 40420;
mem_k_index[8617] = 40422;
mem_k_index[8618] = 40425;
mem_k_index[8619] = 40428;
mem_k_index[8620] = 40430;
mem_k_index[8621] = 40433;
mem_k_index[8622] = 40435;
mem_k_index[8623] = 40438;
mem_k_index[8624] = 40440;
mem_k_index[8625] = 40443;
mem_k_index[8626] = 40445;
mem_k_index[8627] = 40448;
mem_k_index[8628] = 40450;
mem_k_index[8629] = 40453;
mem_k_index[8630] = 40455;
mem_k_index[8631] = 40458;
mem_k_index[8632] = 40460;
mem_k_index[8633] = 40463;
mem_k_index[8634] = 40465;
mem_k_index[8635] = 40468;
mem_k_index[8636] = 40470;
mem_k_index[8637] = 40473;
mem_k_index[8638] = 40475;
mem_k_index[8639] = 40478;
mem_k_index[8640] = 40480;
mem_k_index[8641] = 40483;
mem_k_index[8642] = 40485;
mem_k_index[8643] = 40488;
mem_k_index[8644] = 40490;
mem_k_index[8645] = 40493;
mem_k_index[8646] = 40495;
mem_k_index[8647] = 40498;
mem_k_index[8648] = 40500;
mem_k_index[8649] = 40503;
mem_k_index[8650] = 40505;
mem_k_index[8651] = 40508;
mem_k_index[8652] = 40510;
mem_k_index[8653] = 40513;
mem_k_index[8654] = 40515;
mem_k_index[8655] = 40518;
mem_k_index[8656] = 40520;
mem_k_index[8657] = 40523;
mem_k_index[8658] = 40525;
mem_k_index[8659] = 40528;
mem_k_index[8660] = 40530;
mem_k_index[8661] = 40533;
mem_k_index[8662] = 40536;
mem_k_index[8663] = 40538;
mem_k_index[8664] = 40541;
mem_k_index[8665] = 40543;
mem_k_index[8666] = 40546;
mem_k_index[8667] = 40548;
mem_k_index[8668] = 40551;
mem_k_index[8669] = 40553;
mem_k_index[8670] = 40556;
mem_k_index[8671] = 40558;
mem_k_index[8672] = 40561;
mem_k_index[8673] = 40563;
mem_k_index[8674] = 40566;
mem_k_index[8675] = 40568;
mem_k_index[8676] = 40571;
mem_k_index[8677] = 40573;
mem_k_index[8678] = 40576;
mem_k_index[8679] = 40578;
mem_k_index[8680] = 40581;
mem_k_index[8681] = 40583;
mem_k_index[8682] = 40586;
mem_k_index[8683] = 40588;
mem_k_index[8684] = 40591;
mem_k_index[8685] = 40593;
mem_k_index[8686] = 40596;
mem_k_index[8687] = 40598;
mem_k_index[8688] = 40601;
mem_k_index[8689] = 40603;
mem_k_index[8690] = 40606;
mem_k_index[8691] = 40608;
mem_k_index[8692] = 40611;
mem_k_index[8693] = 40613;
mem_k_index[8694] = 40616;
mem_k_index[8695] = 40618;
mem_k_index[8696] = 40621;
mem_k_index[8697] = 40623;
mem_k_index[8698] = 40626;
mem_k_index[8699] = 40628;
mem_k_index[8700] = 40631;
mem_k_index[8701] = 40633;
mem_k_index[8702] = 40636;
mem_k_index[8703] = 40638;
mem_k_index[8704] = 40640;
mem_k_index[8705] = 40642;
mem_k_index[8706] = 40645;
mem_k_index[8707] = 40647;
mem_k_index[8708] = 40650;
mem_k_index[8709] = 40652;
mem_k_index[8710] = 40655;
mem_k_index[8711] = 40657;
mem_k_index[8712] = 40660;
mem_k_index[8713] = 40662;
mem_k_index[8714] = 40665;
mem_k_index[8715] = 40667;
mem_k_index[8716] = 40670;
mem_k_index[8717] = 40672;
mem_k_index[8718] = 40675;
mem_k_index[8719] = 40677;
mem_k_index[8720] = 40680;
mem_k_index[8721] = 40682;
mem_k_index[8722] = 40685;
mem_k_index[8723] = 40687;
mem_k_index[8724] = 40690;
mem_k_index[8725] = 40692;
mem_k_index[8726] = 40695;
mem_k_index[8727] = 40697;
mem_k_index[8728] = 40700;
mem_k_index[8729] = 40702;
mem_k_index[8730] = 40705;
mem_k_index[8731] = 40707;
mem_k_index[8732] = 40710;
mem_k_index[8733] = 40712;
mem_k_index[8734] = 40715;
mem_k_index[8735] = 40717;
mem_k_index[8736] = 40720;
mem_k_index[8737] = 40722;
mem_k_index[8738] = 40725;
mem_k_index[8739] = 40727;
mem_k_index[8740] = 40730;
mem_k_index[8741] = 40732;
mem_k_index[8742] = 40735;
mem_k_index[8743] = 40737;
mem_k_index[8744] = 40740;
mem_k_index[8745] = 40742;
mem_k_index[8746] = 40745;
mem_k_index[8747] = 40748;
mem_k_index[8748] = 40750;
mem_k_index[8749] = 40753;
mem_k_index[8750] = 40755;
mem_k_index[8751] = 40758;
mem_k_index[8752] = 40760;
mem_k_index[8753] = 40763;
mem_k_index[8754] = 40765;
mem_k_index[8755] = 40768;
mem_k_index[8756] = 40770;
mem_k_index[8757] = 40773;
mem_k_index[8758] = 40775;
mem_k_index[8759] = 40778;
mem_k_index[8760] = 40780;
mem_k_index[8761] = 40783;
mem_k_index[8762] = 40785;
mem_k_index[8763] = 40788;
mem_k_index[8764] = 40790;
mem_k_index[8765] = 40793;
mem_k_index[8766] = 40795;
mem_k_index[8767] = 40798;
mem_k_index[8768] = 40800;
mem_k_index[8769] = 40803;
mem_k_index[8770] = 40805;
mem_k_index[8771] = 40808;
mem_k_index[8772] = 40810;
mem_k_index[8773] = 40813;
mem_k_index[8774] = 40815;
mem_k_index[8775] = 40818;
mem_k_index[8776] = 40820;
mem_k_index[8777] = 40823;
mem_k_index[8778] = 40825;
mem_k_index[8779] = 40828;
mem_k_index[8780] = 40830;
mem_k_index[8781] = 40833;
mem_k_index[8782] = 40835;
mem_k_index[8783] = 40838;
mem_k_index[8784] = 40840;
mem_k_index[8785] = 40843;
mem_k_index[8786] = 40845;
mem_k_index[8787] = 40848;
mem_k_index[8788] = 40850;
mem_k_index[8789] = 40853;
mem_k_index[8790] = 40856;
mem_k_index[8791] = 40858;
mem_k_index[8792] = 40861;
mem_k_index[8793] = 40863;
mem_k_index[8794] = 40866;
mem_k_index[8795] = 40868;
mem_k_index[8796] = 40871;
mem_k_index[8797] = 40873;
mem_k_index[8798] = 40876;
mem_k_index[8799] = 40878;
mem_k_index[8800] = 40881;
mem_k_index[8801] = 40883;
mem_k_index[8802] = 40886;
mem_k_index[8803] = 40888;
mem_k_index[8804] = 40891;
mem_k_index[8805] = 40893;
mem_k_index[8806] = 40896;
mem_k_index[8807] = 40898;
mem_k_index[8808] = 40901;
mem_k_index[8809] = 40903;
mem_k_index[8810] = 40906;
mem_k_index[8811] = 40908;
mem_k_index[8812] = 40911;
mem_k_index[8813] = 40913;
mem_k_index[8814] = 40916;
mem_k_index[8815] = 40918;
mem_k_index[8816] = 40921;
mem_k_index[8817] = 40923;
mem_k_index[8818] = 40926;
mem_k_index[8819] = 40928;
mem_k_index[8820] = 40931;
mem_k_index[8821] = 40933;
mem_k_index[8822] = 40936;
mem_k_index[8823] = 40938;
mem_k_index[8824] = 40941;
mem_k_index[8825] = 40943;
mem_k_index[8826] = 40946;
mem_k_index[8827] = 40948;
mem_k_index[8828] = 40951;
mem_k_index[8829] = 40953;
mem_k_index[8830] = 40956;
mem_k_index[8831] = 40958;
mem_k_index[8832] = 41280;
mem_k_index[8833] = 41282;
mem_k_index[8834] = 41285;
mem_k_index[8835] = 41287;
mem_k_index[8836] = 41290;
mem_k_index[8837] = 41292;
mem_k_index[8838] = 41295;
mem_k_index[8839] = 41297;
mem_k_index[8840] = 41300;
mem_k_index[8841] = 41302;
mem_k_index[8842] = 41305;
mem_k_index[8843] = 41307;
mem_k_index[8844] = 41310;
mem_k_index[8845] = 41312;
mem_k_index[8846] = 41315;
mem_k_index[8847] = 41317;
mem_k_index[8848] = 41320;
mem_k_index[8849] = 41322;
mem_k_index[8850] = 41325;
mem_k_index[8851] = 41327;
mem_k_index[8852] = 41330;
mem_k_index[8853] = 41332;
mem_k_index[8854] = 41335;
mem_k_index[8855] = 41337;
mem_k_index[8856] = 41340;
mem_k_index[8857] = 41342;
mem_k_index[8858] = 41345;
mem_k_index[8859] = 41347;
mem_k_index[8860] = 41350;
mem_k_index[8861] = 41352;
mem_k_index[8862] = 41355;
mem_k_index[8863] = 41357;
mem_k_index[8864] = 41360;
mem_k_index[8865] = 41362;
mem_k_index[8866] = 41365;
mem_k_index[8867] = 41367;
mem_k_index[8868] = 41370;
mem_k_index[8869] = 41372;
mem_k_index[8870] = 41375;
mem_k_index[8871] = 41377;
mem_k_index[8872] = 41380;
mem_k_index[8873] = 41382;
mem_k_index[8874] = 41385;
mem_k_index[8875] = 41388;
mem_k_index[8876] = 41390;
mem_k_index[8877] = 41393;
mem_k_index[8878] = 41395;
mem_k_index[8879] = 41398;
mem_k_index[8880] = 41400;
mem_k_index[8881] = 41403;
mem_k_index[8882] = 41405;
mem_k_index[8883] = 41408;
mem_k_index[8884] = 41410;
mem_k_index[8885] = 41413;
mem_k_index[8886] = 41415;
mem_k_index[8887] = 41418;
mem_k_index[8888] = 41420;
mem_k_index[8889] = 41423;
mem_k_index[8890] = 41425;
mem_k_index[8891] = 41428;
mem_k_index[8892] = 41430;
mem_k_index[8893] = 41433;
mem_k_index[8894] = 41435;
mem_k_index[8895] = 41438;
mem_k_index[8896] = 41440;
mem_k_index[8897] = 41443;
mem_k_index[8898] = 41445;
mem_k_index[8899] = 41448;
mem_k_index[8900] = 41450;
mem_k_index[8901] = 41453;
mem_k_index[8902] = 41455;
mem_k_index[8903] = 41458;
mem_k_index[8904] = 41460;
mem_k_index[8905] = 41463;
mem_k_index[8906] = 41465;
mem_k_index[8907] = 41468;
mem_k_index[8908] = 41470;
mem_k_index[8909] = 41473;
mem_k_index[8910] = 41475;
mem_k_index[8911] = 41478;
mem_k_index[8912] = 41480;
mem_k_index[8913] = 41483;
mem_k_index[8914] = 41485;
mem_k_index[8915] = 41488;
mem_k_index[8916] = 41490;
mem_k_index[8917] = 41493;
mem_k_index[8918] = 41496;
mem_k_index[8919] = 41498;
mem_k_index[8920] = 41501;
mem_k_index[8921] = 41503;
mem_k_index[8922] = 41506;
mem_k_index[8923] = 41508;
mem_k_index[8924] = 41511;
mem_k_index[8925] = 41513;
mem_k_index[8926] = 41516;
mem_k_index[8927] = 41518;
mem_k_index[8928] = 41521;
mem_k_index[8929] = 41523;
mem_k_index[8930] = 41526;
mem_k_index[8931] = 41528;
mem_k_index[8932] = 41531;
mem_k_index[8933] = 41533;
mem_k_index[8934] = 41536;
mem_k_index[8935] = 41538;
mem_k_index[8936] = 41541;
mem_k_index[8937] = 41543;
mem_k_index[8938] = 41546;
mem_k_index[8939] = 41548;
mem_k_index[8940] = 41551;
mem_k_index[8941] = 41553;
mem_k_index[8942] = 41556;
mem_k_index[8943] = 41558;
mem_k_index[8944] = 41561;
mem_k_index[8945] = 41563;
mem_k_index[8946] = 41566;
mem_k_index[8947] = 41568;
mem_k_index[8948] = 41571;
mem_k_index[8949] = 41573;
mem_k_index[8950] = 41576;
mem_k_index[8951] = 41578;
mem_k_index[8952] = 41581;
mem_k_index[8953] = 41583;
mem_k_index[8954] = 41586;
mem_k_index[8955] = 41588;
mem_k_index[8956] = 41591;
mem_k_index[8957] = 41593;
mem_k_index[8958] = 41596;
mem_k_index[8959] = 41598;
mem_k_index[8960] = 41920;
mem_k_index[8961] = 41922;
mem_k_index[8962] = 41925;
mem_k_index[8963] = 41927;
mem_k_index[8964] = 41930;
mem_k_index[8965] = 41932;
mem_k_index[8966] = 41935;
mem_k_index[8967] = 41937;
mem_k_index[8968] = 41940;
mem_k_index[8969] = 41942;
mem_k_index[8970] = 41945;
mem_k_index[8971] = 41947;
mem_k_index[8972] = 41950;
mem_k_index[8973] = 41952;
mem_k_index[8974] = 41955;
mem_k_index[8975] = 41957;
mem_k_index[8976] = 41960;
mem_k_index[8977] = 41962;
mem_k_index[8978] = 41965;
mem_k_index[8979] = 41967;
mem_k_index[8980] = 41970;
mem_k_index[8981] = 41972;
mem_k_index[8982] = 41975;
mem_k_index[8983] = 41977;
mem_k_index[8984] = 41980;
mem_k_index[8985] = 41982;
mem_k_index[8986] = 41985;
mem_k_index[8987] = 41987;
mem_k_index[8988] = 41990;
mem_k_index[8989] = 41992;
mem_k_index[8990] = 41995;
mem_k_index[8991] = 41997;
mem_k_index[8992] = 42000;
mem_k_index[8993] = 42002;
mem_k_index[8994] = 42005;
mem_k_index[8995] = 42007;
mem_k_index[8996] = 42010;
mem_k_index[8997] = 42012;
mem_k_index[8998] = 42015;
mem_k_index[8999] = 42017;
mem_k_index[9000] = 42020;
mem_k_index[9001] = 42022;
mem_k_index[9002] = 42025;
mem_k_index[9003] = 42028;
mem_k_index[9004] = 42030;
mem_k_index[9005] = 42033;
mem_k_index[9006] = 42035;
mem_k_index[9007] = 42038;
mem_k_index[9008] = 42040;
mem_k_index[9009] = 42043;
mem_k_index[9010] = 42045;
mem_k_index[9011] = 42048;
mem_k_index[9012] = 42050;
mem_k_index[9013] = 42053;
mem_k_index[9014] = 42055;
mem_k_index[9015] = 42058;
mem_k_index[9016] = 42060;
mem_k_index[9017] = 42063;
mem_k_index[9018] = 42065;
mem_k_index[9019] = 42068;
mem_k_index[9020] = 42070;
mem_k_index[9021] = 42073;
mem_k_index[9022] = 42075;
mem_k_index[9023] = 42078;
mem_k_index[9024] = 42080;
mem_k_index[9025] = 42083;
mem_k_index[9026] = 42085;
mem_k_index[9027] = 42088;
mem_k_index[9028] = 42090;
mem_k_index[9029] = 42093;
mem_k_index[9030] = 42095;
mem_k_index[9031] = 42098;
mem_k_index[9032] = 42100;
mem_k_index[9033] = 42103;
mem_k_index[9034] = 42105;
mem_k_index[9035] = 42108;
mem_k_index[9036] = 42110;
mem_k_index[9037] = 42113;
mem_k_index[9038] = 42115;
mem_k_index[9039] = 42118;
mem_k_index[9040] = 42120;
mem_k_index[9041] = 42123;
mem_k_index[9042] = 42125;
mem_k_index[9043] = 42128;
mem_k_index[9044] = 42130;
mem_k_index[9045] = 42133;
mem_k_index[9046] = 42136;
mem_k_index[9047] = 42138;
mem_k_index[9048] = 42141;
mem_k_index[9049] = 42143;
mem_k_index[9050] = 42146;
mem_k_index[9051] = 42148;
mem_k_index[9052] = 42151;
mem_k_index[9053] = 42153;
mem_k_index[9054] = 42156;
mem_k_index[9055] = 42158;
mem_k_index[9056] = 42161;
mem_k_index[9057] = 42163;
mem_k_index[9058] = 42166;
mem_k_index[9059] = 42168;
mem_k_index[9060] = 42171;
mem_k_index[9061] = 42173;
mem_k_index[9062] = 42176;
mem_k_index[9063] = 42178;
mem_k_index[9064] = 42181;
mem_k_index[9065] = 42183;
mem_k_index[9066] = 42186;
mem_k_index[9067] = 42188;
mem_k_index[9068] = 42191;
mem_k_index[9069] = 42193;
mem_k_index[9070] = 42196;
mem_k_index[9071] = 42198;
mem_k_index[9072] = 42201;
mem_k_index[9073] = 42203;
mem_k_index[9074] = 42206;
mem_k_index[9075] = 42208;
mem_k_index[9076] = 42211;
mem_k_index[9077] = 42213;
mem_k_index[9078] = 42216;
mem_k_index[9079] = 42218;
mem_k_index[9080] = 42221;
mem_k_index[9081] = 42223;
mem_k_index[9082] = 42226;
mem_k_index[9083] = 42228;
mem_k_index[9084] = 42231;
mem_k_index[9085] = 42233;
mem_k_index[9086] = 42236;
mem_k_index[9087] = 42238;
mem_k_index[9088] = 42560;
mem_k_index[9089] = 42562;
mem_k_index[9090] = 42565;
mem_k_index[9091] = 42567;
mem_k_index[9092] = 42570;
mem_k_index[9093] = 42572;
mem_k_index[9094] = 42575;
mem_k_index[9095] = 42577;
mem_k_index[9096] = 42580;
mem_k_index[9097] = 42582;
mem_k_index[9098] = 42585;
mem_k_index[9099] = 42587;
mem_k_index[9100] = 42590;
mem_k_index[9101] = 42592;
mem_k_index[9102] = 42595;
mem_k_index[9103] = 42597;
mem_k_index[9104] = 42600;
mem_k_index[9105] = 42602;
mem_k_index[9106] = 42605;
mem_k_index[9107] = 42607;
mem_k_index[9108] = 42610;
mem_k_index[9109] = 42612;
mem_k_index[9110] = 42615;
mem_k_index[9111] = 42617;
mem_k_index[9112] = 42620;
mem_k_index[9113] = 42622;
mem_k_index[9114] = 42625;
mem_k_index[9115] = 42627;
mem_k_index[9116] = 42630;
mem_k_index[9117] = 42632;
mem_k_index[9118] = 42635;
mem_k_index[9119] = 42637;
mem_k_index[9120] = 42640;
mem_k_index[9121] = 42642;
mem_k_index[9122] = 42645;
mem_k_index[9123] = 42647;
mem_k_index[9124] = 42650;
mem_k_index[9125] = 42652;
mem_k_index[9126] = 42655;
mem_k_index[9127] = 42657;
mem_k_index[9128] = 42660;
mem_k_index[9129] = 42662;
mem_k_index[9130] = 42665;
mem_k_index[9131] = 42668;
mem_k_index[9132] = 42670;
mem_k_index[9133] = 42673;
mem_k_index[9134] = 42675;
mem_k_index[9135] = 42678;
mem_k_index[9136] = 42680;
mem_k_index[9137] = 42683;
mem_k_index[9138] = 42685;
mem_k_index[9139] = 42688;
mem_k_index[9140] = 42690;
mem_k_index[9141] = 42693;
mem_k_index[9142] = 42695;
mem_k_index[9143] = 42698;
mem_k_index[9144] = 42700;
mem_k_index[9145] = 42703;
mem_k_index[9146] = 42705;
mem_k_index[9147] = 42708;
mem_k_index[9148] = 42710;
mem_k_index[9149] = 42713;
mem_k_index[9150] = 42715;
mem_k_index[9151] = 42718;
mem_k_index[9152] = 42720;
mem_k_index[9153] = 42723;
mem_k_index[9154] = 42725;
mem_k_index[9155] = 42728;
mem_k_index[9156] = 42730;
mem_k_index[9157] = 42733;
mem_k_index[9158] = 42735;
mem_k_index[9159] = 42738;
mem_k_index[9160] = 42740;
mem_k_index[9161] = 42743;
mem_k_index[9162] = 42745;
mem_k_index[9163] = 42748;
mem_k_index[9164] = 42750;
mem_k_index[9165] = 42753;
mem_k_index[9166] = 42755;
mem_k_index[9167] = 42758;
mem_k_index[9168] = 42760;
mem_k_index[9169] = 42763;
mem_k_index[9170] = 42765;
mem_k_index[9171] = 42768;
mem_k_index[9172] = 42770;
mem_k_index[9173] = 42773;
mem_k_index[9174] = 42776;
mem_k_index[9175] = 42778;
mem_k_index[9176] = 42781;
mem_k_index[9177] = 42783;
mem_k_index[9178] = 42786;
mem_k_index[9179] = 42788;
mem_k_index[9180] = 42791;
mem_k_index[9181] = 42793;
mem_k_index[9182] = 42796;
mem_k_index[9183] = 42798;
mem_k_index[9184] = 42801;
mem_k_index[9185] = 42803;
mem_k_index[9186] = 42806;
mem_k_index[9187] = 42808;
mem_k_index[9188] = 42811;
mem_k_index[9189] = 42813;
mem_k_index[9190] = 42816;
mem_k_index[9191] = 42818;
mem_k_index[9192] = 42821;
mem_k_index[9193] = 42823;
mem_k_index[9194] = 42826;
mem_k_index[9195] = 42828;
mem_k_index[9196] = 42831;
mem_k_index[9197] = 42833;
mem_k_index[9198] = 42836;
mem_k_index[9199] = 42838;
mem_k_index[9200] = 42841;
mem_k_index[9201] = 42843;
mem_k_index[9202] = 42846;
mem_k_index[9203] = 42848;
mem_k_index[9204] = 42851;
mem_k_index[9205] = 42853;
mem_k_index[9206] = 42856;
mem_k_index[9207] = 42858;
mem_k_index[9208] = 42861;
mem_k_index[9209] = 42863;
mem_k_index[9210] = 42866;
mem_k_index[9211] = 42868;
mem_k_index[9212] = 42871;
mem_k_index[9213] = 42873;
mem_k_index[9214] = 42876;
mem_k_index[9215] = 42878;
mem_k_index[9216] = 43200;
mem_k_index[9217] = 43202;
mem_k_index[9218] = 43205;
mem_k_index[9219] = 43207;
mem_k_index[9220] = 43210;
mem_k_index[9221] = 43212;
mem_k_index[9222] = 43215;
mem_k_index[9223] = 43217;
mem_k_index[9224] = 43220;
mem_k_index[9225] = 43222;
mem_k_index[9226] = 43225;
mem_k_index[9227] = 43227;
mem_k_index[9228] = 43230;
mem_k_index[9229] = 43232;
mem_k_index[9230] = 43235;
mem_k_index[9231] = 43237;
mem_k_index[9232] = 43240;
mem_k_index[9233] = 43242;
mem_k_index[9234] = 43245;
mem_k_index[9235] = 43247;
mem_k_index[9236] = 43250;
mem_k_index[9237] = 43252;
mem_k_index[9238] = 43255;
mem_k_index[9239] = 43257;
mem_k_index[9240] = 43260;
mem_k_index[9241] = 43262;
mem_k_index[9242] = 43265;
mem_k_index[9243] = 43267;
mem_k_index[9244] = 43270;
mem_k_index[9245] = 43272;
mem_k_index[9246] = 43275;
mem_k_index[9247] = 43277;
mem_k_index[9248] = 43280;
mem_k_index[9249] = 43282;
mem_k_index[9250] = 43285;
mem_k_index[9251] = 43287;
mem_k_index[9252] = 43290;
mem_k_index[9253] = 43292;
mem_k_index[9254] = 43295;
mem_k_index[9255] = 43297;
mem_k_index[9256] = 43300;
mem_k_index[9257] = 43302;
mem_k_index[9258] = 43305;
mem_k_index[9259] = 43308;
mem_k_index[9260] = 43310;
mem_k_index[9261] = 43313;
mem_k_index[9262] = 43315;
mem_k_index[9263] = 43318;
mem_k_index[9264] = 43320;
mem_k_index[9265] = 43323;
mem_k_index[9266] = 43325;
mem_k_index[9267] = 43328;
mem_k_index[9268] = 43330;
mem_k_index[9269] = 43333;
mem_k_index[9270] = 43335;
mem_k_index[9271] = 43338;
mem_k_index[9272] = 43340;
mem_k_index[9273] = 43343;
mem_k_index[9274] = 43345;
mem_k_index[9275] = 43348;
mem_k_index[9276] = 43350;
mem_k_index[9277] = 43353;
mem_k_index[9278] = 43355;
mem_k_index[9279] = 43358;
mem_k_index[9280] = 43360;
mem_k_index[9281] = 43363;
mem_k_index[9282] = 43365;
mem_k_index[9283] = 43368;
mem_k_index[9284] = 43370;
mem_k_index[9285] = 43373;
mem_k_index[9286] = 43375;
mem_k_index[9287] = 43378;
mem_k_index[9288] = 43380;
mem_k_index[9289] = 43383;
mem_k_index[9290] = 43385;
mem_k_index[9291] = 43388;
mem_k_index[9292] = 43390;
mem_k_index[9293] = 43393;
mem_k_index[9294] = 43395;
mem_k_index[9295] = 43398;
mem_k_index[9296] = 43400;
mem_k_index[9297] = 43403;
mem_k_index[9298] = 43405;
mem_k_index[9299] = 43408;
mem_k_index[9300] = 43410;
mem_k_index[9301] = 43413;
mem_k_index[9302] = 43416;
mem_k_index[9303] = 43418;
mem_k_index[9304] = 43421;
mem_k_index[9305] = 43423;
mem_k_index[9306] = 43426;
mem_k_index[9307] = 43428;
mem_k_index[9308] = 43431;
mem_k_index[9309] = 43433;
mem_k_index[9310] = 43436;
mem_k_index[9311] = 43438;
mem_k_index[9312] = 43441;
mem_k_index[9313] = 43443;
mem_k_index[9314] = 43446;
mem_k_index[9315] = 43448;
mem_k_index[9316] = 43451;
mem_k_index[9317] = 43453;
mem_k_index[9318] = 43456;
mem_k_index[9319] = 43458;
mem_k_index[9320] = 43461;
mem_k_index[9321] = 43463;
mem_k_index[9322] = 43466;
mem_k_index[9323] = 43468;
mem_k_index[9324] = 43471;
mem_k_index[9325] = 43473;
mem_k_index[9326] = 43476;
mem_k_index[9327] = 43478;
mem_k_index[9328] = 43481;
mem_k_index[9329] = 43483;
mem_k_index[9330] = 43486;
mem_k_index[9331] = 43488;
mem_k_index[9332] = 43491;
mem_k_index[9333] = 43493;
mem_k_index[9334] = 43496;
mem_k_index[9335] = 43498;
mem_k_index[9336] = 43501;
mem_k_index[9337] = 43503;
mem_k_index[9338] = 43506;
mem_k_index[9339] = 43508;
mem_k_index[9340] = 43511;
mem_k_index[9341] = 43513;
mem_k_index[9342] = 43516;
mem_k_index[9343] = 43518;
mem_k_index[9344] = 43840;
mem_k_index[9345] = 43842;
mem_k_index[9346] = 43845;
mem_k_index[9347] = 43847;
mem_k_index[9348] = 43850;
mem_k_index[9349] = 43852;
mem_k_index[9350] = 43855;
mem_k_index[9351] = 43857;
mem_k_index[9352] = 43860;
mem_k_index[9353] = 43862;
mem_k_index[9354] = 43865;
mem_k_index[9355] = 43867;
mem_k_index[9356] = 43870;
mem_k_index[9357] = 43872;
mem_k_index[9358] = 43875;
mem_k_index[9359] = 43877;
mem_k_index[9360] = 43880;
mem_k_index[9361] = 43882;
mem_k_index[9362] = 43885;
mem_k_index[9363] = 43887;
mem_k_index[9364] = 43890;
mem_k_index[9365] = 43892;
mem_k_index[9366] = 43895;
mem_k_index[9367] = 43897;
mem_k_index[9368] = 43900;
mem_k_index[9369] = 43902;
mem_k_index[9370] = 43905;
mem_k_index[9371] = 43907;
mem_k_index[9372] = 43910;
mem_k_index[9373] = 43912;
mem_k_index[9374] = 43915;
mem_k_index[9375] = 43917;
mem_k_index[9376] = 43920;
mem_k_index[9377] = 43922;
mem_k_index[9378] = 43925;
mem_k_index[9379] = 43927;
mem_k_index[9380] = 43930;
mem_k_index[9381] = 43932;
mem_k_index[9382] = 43935;
mem_k_index[9383] = 43937;
mem_k_index[9384] = 43940;
mem_k_index[9385] = 43942;
mem_k_index[9386] = 43945;
mem_k_index[9387] = 43948;
mem_k_index[9388] = 43950;
mem_k_index[9389] = 43953;
mem_k_index[9390] = 43955;
mem_k_index[9391] = 43958;
mem_k_index[9392] = 43960;
mem_k_index[9393] = 43963;
mem_k_index[9394] = 43965;
mem_k_index[9395] = 43968;
mem_k_index[9396] = 43970;
mem_k_index[9397] = 43973;
mem_k_index[9398] = 43975;
mem_k_index[9399] = 43978;
mem_k_index[9400] = 43980;
mem_k_index[9401] = 43983;
mem_k_index[9402] = 43985;
mem_k_index[9403] = 43988;
mem_k_index[9404] = 43990;
mem_k_index[9405] = 43993;
mem_k_index[9406] = 43995;
mem_k_index[9407] = 43998;
mem_k_index[9408] = 44000;
mem_k_index[9409] = 44003;
mem_k_index[9410] = 44005;
mem_k_index[9411] = 44008;
mem_k_index[9412] = 44010;
mem_k_index[9413] = 44013;
mem_k_index[9414] = 44015;
mem_k_index[9415] = 44018;
mem_k_index[9416] = 44020;
mem_k_index[9417] = 44023;
mem_k_index[9418] = 44025;
mem_k_index[9419] = 44028;
mem_k_index[9420] = 44030;
mem_k_index[9421] = 44033;
mem_k_index[9422] = 44035;
mem_k_index[9423] = 44038;
mem_k_index[9424] = 44040;
mem_k_index[9425] = 44043;
mem_k_index[9426] = 44045;
mem_k_index[9427] = 44048;
mem_k_index[9428] = 44050;
mem_k_index[9429] = 44053;
mem_k_index[9430] = 44056;
mem_k_index[9431] = 44058;
mem_k_index[9432] = 44061;
mem_k_index[9433] = 44063;
mem_k_index[9434] = 44066;
mem_k_index[9435] = 44068;
mem_k_index[9436] = 44071;
mem_k_index[9437] = 44073;
mem_k_index[9438] = 44076;
mem_k_index[9439] = 44078;
mem_k_index[9440] = 44081;
mem_k_index[9441] = 44083;
mem_k_index[9442] = 44086;
mem_k_index[9443] = 44088;
mem_k_index[9444] = 44091;
mem_k_index[9445] = 44093;
mem_k_index[9446] = 44096;
mem_k_index[9447] = 44098;
mem_k_index[9448] = 44101;
mem_k_index[9449] = 44103;
mem_k_index[9450] = 44106;
mem_k_index[9451] = 44108;
mem_k_index[9452] = 44111;
mem_k_index[9453] = 44113;
mem_k_index[9454] = 44116;
mem_k_index[9455] = 44118;
mem_k_index[9456] = 44121;
mem_k_index[9457] = 44123;
mem_k_index[9458] = 44126;
mem_k_index[9459] = 44128;
mem_k_index[9460] = 44131;
mem_k_index[9461] = 44133;
mem_k_index[9462] = 44136;
mem_k_index[9463] = 44138;
mem_k_index[9464] = 44141;
mem_k_index[9465] = 44143;
mem_k_index[9466] = 44146;
mem_k_index[9467] = 44148;
mem_k_index[9468] = 44151;
mem_k_index[9469] = 44153;
mem_k_index[9470] = 44156;
mem_k_index[9471] = 44158;
mem_k_index[9472] = 44480;
mem_k_index[9473] = 44482;
mem_k_index[9474] = 44485;
mem_k_index[9475] = 44487;
mem_k_index[9476] = 44490;
mem_k_index[9477] = 44492;
mem_k_index[9478] = 44495;
mem_k_index[9479] = 44497;
mem_k_index[9480] = 44500;
mem_k_index[9481] = 44502;
mem_k_index[9482] = 44505;
mem_k_index[9483] = 44507;
mem_k_index[9484] = 44510;
mem_k_index[9485] = 44512;
mem_k_index[9486] = 44515;
mem_k_index[9487] = 44517;
mem_k_index[9488] = 44520;
mem_k_index[9489] = 44522;
mem_k_index[9490] = 44525;
mem_k_index[9491] = 44527;
mem_k_index[9492] = 44530;
mem_k_index[9493] = 44532;
mem_k_index[9494] = 44535;
mem_k_index[9495] = 44537;
mem_k_index[9496] = 44540;
mem_k_index[9497] = 44542;
mem_k_index[9498] = 44545;
mem_k_index[9499] = 44547;
mem_k_index[9500] = 44550;
mem_k_index[9501] = 44552;
mem_k_index[9502] = 44555;
mem_k_index[9503] = 44557;
mem_k_index[9504] = 44560;
mem_k_index[9505] = 44562;
mem_k_index[9506] = 44565;
mem_k_index[9507] = 44567;
mem_k_index[9508] = 44570;
mem_k_index[9509] = 44572;
mem_k_index[9510] = 44575;
mem_k_index[9511] = 44577;
mem_k_index[9512] = 44580;
mem_k_index[9513] = 44582;
mem_k_index[9514] = 44585;
mem_k_index[9515] = 44588;
mem_k_index[9516] = 44590;
mem_k_index[9517] = 44593;
mem_k_index[9518] = 44595;
mem_k_index[9519] = 44598;
mem_k_index[9520] = 44600;
mem_k_index[9521] = 44603;
mem_k_index[9522] = 44605;
mem_k_index[9523] = 44608;
mem_k_index[9524] = 44610;
mem_k_index[9525] = 44613;
mem_k_index[9526] = 44615;
mem_k_index[9527] = 44618;
mem_k_index[9528] = 44620;
mem_k_index[9529] = 44623;
mem_k_index[9530] = 44625;
mem_k_index[9531] = 44628;
mem_k_index[9532] = 44630;
mem_k_index[9533] = 44633;
mem_k_index[9534] = 44635;
mem_k_index[9535] = 44638;
mem_k_index[9536] = 44640;
mem_k_index[9537] = 44643;
mem_k_index[9538] = 44645;
mem_k_index[9539] = 44648;
mem_k_index[9540] = 44650;
mem_k_index[9541] = 44653;
mem_k_index[9542] = 44655;
mem_k_index[9543] = 44658;
mem_k_index[9544] = 44660;
mem_k_index[9545] = 44663;
mem_k_index[9546] = 44665;
mem_k_index[9547] = 44668;
mem_k_index[9548] = 44670;
mem_k_index[9549] = 44673;
mem_k_index[9550] = 44675;
mem_k_index[9551] = 44678;
mem_k_index[9552] = 44680;
mem_k_index[9553] = 44683;
mem_k_index[9554] = 44685;
mem_k_index[9555] = 44688;
mem_k_index[9556] = 44690;
mem_k_index[9557] = 44693;
mem_k_index[9558] = 44696;
mem_k_index[9559] = 44698;
mem_k_index[9560] = 44701;
mem_k_index[9561] = 44703;
mem_k_index[9562] = 44706;
mem_k_index[9563] = 44708;
mem_k_index[9564] = 44711;
mem_k_index[9565] = 44713;
mem_k_index[9566] = 44716;
mem_k_index[9567] = 44718;
mem_k_index[9568] = 44721;
mem_k_index[9569] = 44723;
mem_k_index[9570] = 44726;
mem_k_index[9571] = 44728;
mem_k_index[9572] = 44731;
mem_k_index[9573] = 44733;
mem_k_index[9574] = 44736;
mem_k_index[9575] = 44738;
mem_k_index[9576] = 44741;
mem_k_index[9577] = 44743;
mem_k_index[9578] = 44746;
mem_k_index[9579] = 44748;
mem_k_index[9580] = 44751;
mem_k_index[9581] = 44753;
mem_k_index[9582] = 44756;
mem_k_index[9583] = 44758;
mem_k_index[9584] = 44761;
mem_k_index[9585] = 44763;
mem_k_index[9586] = 44766;
mem_k_index[9587] = 44768;
mem_k_index[9588] = 44771;
mem_k_index[9589] = 44773;
mem_k_index[9590] = 44776;
mem_k_index[9591] = 44778;
mem_k_index[9592] = 44781;
mem_k_index[9593] = 44783;
mem_k_index[9594] = 44786;
mem_k_index[9595] = 44788;
mem_k_index[9596] = 44791;
mem_k_index[9597] = 44793;
mem_k_index[9598] = 44796;
mem_k_index[9599] = 44798;
mem_k_index[9600] = 45120;
mem_k_index[9601] = 45122;
mem_k_index[9602] = 45125;
mem_k_index[9603] = 45127;
mem_k_index[9604] = 45130;
mem_k_index[9605] = 45132;
mem_k_index[9606] = 45135;
mem_k_index[9607] = 45137;
mem_k_index[9608] = 45140;
mem_k_index[9609] = 45142;
mem_k_index[9610] = 45145;
mem_k_index[9611] = 45147;
mem_k_index[9612] = 45150;
mem_k_index[9613] = 45152;
mem_k_index[9614] = 45155;
mem_k_index[9615] = 45157;
mem_k_index[9616] = 45160;
mem_k_index[9617] = 45162;
mem_k_index[9618] = 45165;
mem_k_index[9619] = 45167;
mem_k_index[9620] = 45170;
mem_k_index[9621] = 45172;
mem_k_index[9622] = 45175;
mem_k_index[9623] = 45177;
mem_k_index[9624] = 45180;
mem_k_index[9625] = 45182;
mem_k_index[9626] = 45185;
mem_k_index[9627] = 45187;
mem_k_index[9628] = 45190;
mem_k_index[9629] = 45192;
mem_k_index[9630] = 45195;
mem_k_index[9631] = 45197;
mem_k_index[9632] = 45200;
mem_k_index[9633] = 45202;
mem_k_index[9634] = 45205;
mem_k_index[9635] = 45207;
mem_k_index[9636] = 45210;
mem_k_index[9637] = 45212;
mem_k_index[9638] = 45215;
mem_k_index[9639] = 45217;
mem_k_index[9640] = 45220;
mem_k_index[9641] = 45222;
mem_k_index[9642] = 45225;
mem_k_index[9643] = 45228;
mem_k_index[9644] = 45230;
mem_k_index[9645] = 45233;
mem_k_index[9646] = 45235;
mem_k_index[9647] = 45238;
mem_k_index[9648] = 45240;
mem_k_index[9649] = 45243;
mem_k_index[9650] = 45245;
mem_k_index[9651] = 45248;
mem_k_index[9652] = 45250;
mem_k_index[9653] = 45253;
mem_k_index[9654] = 45255;
mem_k_index[9655] = 45258;
mem_k_index[9656] = 45260;
mem_k_index[9657] = 45263;
mem_k_index[9658] = 45265;
mem_k_index[9659] = 45268;
mem_k_index[9660] = 45270;
mem_k_index[9661] = 45273;
mem_k_index[9662] = 45275;
mem_k_index[9663] = 45278;
mem_k_index[9664] = 45280;
mem_k_index[9665] = 45283;
mem_k_index[9666] = 45285;
mem_k_index[9667] = 45288;
mem_k_index[9668] = 45290;
mem_k_index[9669] = 45293;
mem_k_index[9670] = 45295;
mem_k_index[9671] = 45298;
mem_k_index[9672] = 45300;
mem_k_index[9673] = 45303;
mem_k_index[9674] = 45305;
mem_k_index[9675] = 45308;
mem_k_index[9676] = 45310;
mem_k_index[9677] = 45313;
mem_k_index[9678] = 45315;
mem_k_index[9679] = 45318;
mem_k_index[9680] = 45320;
mem_k_index[9681] = 45323;
mem_k_index[9682] = 45325;
mem_k_index[9683] = 45328;
mem_k_index[9684] = 45330;
mem_k_index[9685] = 45333;
mem_k_index[9686] = 45336;
mem_k_index[9687] = 45338;
mem_k_index[9688] = 45341;
mem_k_index[9689] = 45343;
mem_k_index[9690] = 45346;
mem_k_index[9691] = 45348;
mem_k_index[9692] = 45351;
mem_k_index[9693] = 45353;
mem_k_index[9694] = 45356;
mem_k_index[9695] = 45358;
mem_k_index[9696] = 45361;
mem_k_index[9697] = 45363;
mem_k_index[9698] = 45366;
mem_k_index[9699] = 45368;
mem_k_index[9700] = 45371;
mem_k_index[9701] = 45373;
mem_k_index[9702] = 45376;
mem_k_index[9703] = 45378;
mem_k_index[9704] = 45381;
mem_k_index[9705] = 45383;
mem_k_index[9706] = 45386;
mem_k_index[9707] = 45388;
mem_k_index[9708] = 45391;
mem_k_index[9709] = 45393;
mem_k_index[9710] = 45396;
mem_k_index[9711] = 45398;
mem_k_index[9712] = 45401;
mem_k_index[9713] = 45403;
mem_k_index[9714] = 45406;
mem_k_index[9715] = 45408;
mem_k_index[9716] = 45411;
mem_k_index[9717] = 45413;
mem_k_index[9718] = 45416;
mem_k_index[9719] = 45418;
mem_k_index[9720] = 45421;
mem_k_index[9721] = 45423;
mem_k_index[9722] = 45426;
mem_k_index[9723] = 45428;
mem_k_index[9724] = 45431;
mem_k_index[9725] = 45433;
mem_k_index[9726] = 45436;
mem_k_index[9727] = 45438;
mem_k_index[9728] = 45760;
mem_k_index[9729] = 45762;
mem_k_index[9730] = 45765;
mem_k_index[9731] = 45767;
mem_k_index[9732] = 45770;
mem_k_index[9733] = 45772;
mem_k_index[9734] = 45775;
mem_k_index[9735] = 45777;
mem_k_index[9736] = 45780;
mem_k_index[9737] = 45782;
mem_k_index[9738] = 45785;
mem_k_index[9739] = 45787;
mem_k_index[9740] = 45790;
mem_k_index[9741] = 45792;
mem_k_index[9742] = 45795;
mem_k_index[9743] = 45797;
mem_k_index[9744] = 45800;
mem_k_index[9745] = 45802;
mem_k_index[9746] = 45805;
mem_k_index[9747] = 45807;
mem_k_index[9748] = 45810;
mem_k_index[9749] = 45812;
mem_k_index[9750] = 45815;
mem_k_index[9751] = 45817;
mem_k_index[9752] = 45820;
mem_k_index[9753] = 45822;
mem_k_index[9754] = 45825;
mem_k_index[9755] = 45827;
mem_k_index[9756] = 45830;
mem_k_index[9757] = 45832;
mem_k_index[9758] = 45835;
mem_k_index[9759] = 45837;
mem_k_index[9760] = 45840;
mem_k_index[9761] = 45842;
mem_k_index[9762] = 45845;
mem_k_index[9763] = 45847;
mem_k_index[9764] = 45850;
mem_k_index[9765] = 45852;
mem_k_index[9766] = 45855;
mem_k_index[9767] = 45857;
mem_k_index[9768] = 45860;
mem_k_index[9769] = 45862;
mem_k_index[9770] = 45865;
mem_k_index[9771] = 45868;
mem_k_index[9772] = 45870;
mem_k_index[9773] = 45873;
mem_k_index[9774] = 45875;
mem_k_index[9775] = 45878;
mem_k_index[9776] = 45880;
mem_k_index[9777] = 45883;
mem_k_index[9778] = 45885;
mem_k_index[9779] = 45888;
mem_k_index[9780] = 45890;
mem_k_index[9781] = 45893;
mem_k_index[9782] = 45895;
mem_k_index[9783] = 45898;
mem_k_index[9784] = 45900;
mem_k_index[9785] = 45903;
mem_k_index[9786] = 45905;
mem_k_index[9787] = 45908;
mem_k_index[9788] = 45910;
mem_k_index[9789] = 45913;
mem_k_index[9790] = 45915;
mem_k_index[9791] = 45918;
mem_k_index[9792] = 45920;
mem_k_index[9793] = 45923;
mem_k_index[9794] = 45925;
mem_k_index[9795] = 45928;
mem_k_index[9796] = 45930;
mem_k_index[9797] = 45933;
mem_k_index[9798] = 45935;
mem_k_index[9799] = 45938;
mem_k_index[9800] = 45940;
mem_k_index[9801] = 45943;
mem_k_index[9802] = 45945;
mem_k_index[9803] = 45948;
mem_k_index[9804] = 45950;
mem_k_index[9805] = 45953;
mem_k_index[9806] = 45955;
mem_k_index[9807] = 45958;
mem_k_index[9808] = 45960;
mem_k_index[9809] = 45963;
mem_k_index[9810] = 45965;
mem_k_index[9811] = 45968;
mem_k_index[9812] = 45970;
mem_k_index[9813] = 45973;
mem_k_index[9814] = 45976;
mem_k_index[9815] = 45978;
mem_k_index[9816] = 45981;
mem_k_index[9817] = 45983;
mem_k_index[9818] = 45986;
mem_k_index[9819] = 45988;
mem_k_index[9820] = 45991;
mem_k_index[9821] = 45993;
mem_k_index[9822] = 45996;
mem_k_index[9823] = 45998;
mem_k_index[9824] = 46001;
mem_k_index[9825] = 46003;
mem_k_index[9826] = 46006;
mem_k_index[9827] = 46008;
mem_k_index[9828] = 46011;
mem_k_index[9829] = 46013;
mem_k_index[9830] = 46016;
mem_k_index[9831] = 46018;
mem_k_index[9832] = 46021;
mem_k_index[9833] = 46023;
mem_k_index[9834] = 46026;
mem_k_index[9835] = 46028;
mem_k_index[9836] = 46031;
mem_k_index[9837] = 46033;
mem_k_index[9838] = 46036;
mem_k_index[9839] = 46038;
mem_k_index[9840] = 46041;
mem_k_index[9841] = 46043;
mem_k_index[9842] = 46046;
mem_k_index[9843] = 46048;
mem_k_index[9844] = 46051;
mem_k_index[9845] = 46053;
mem_k_index[9846] = 46056;
mem_k_index[9847] = 46058;
mem_k_index[9848] = 46061;
mem_k_index[9849] = 46063;
mem_k_index[9850] = 46066;
mem_k_index[9851] = 46068;
mem_k_index[9852] = 46071;
mem_k_index[9853] = 46073;
mem_k_index[9854] = 46076;
mem_k_index[9855] = 46078;
mem_k_index[9856] = 46080;
mem_k_index[9857] = 46082;
mem_k_index[9858] = 46085;
mem_k_index[9859] = 46087;
mem_k_index[9860] = 46090;
mem_k_index[9861] = 46092;
mem_k_index[9862] = 46095;
mem_k_index[9863] = 46097;
mem_k_index[9864] = 46100;
mem_k_index[9865] = 46102;
mem_k_index[9866] = 46105;
mem_k_index[9867] = 46107;
mem_k_index[9868] = 46110;
mem_k_index[9869] = 46112;
mem_k_index[9870] = 46115;
mem_k_index[9871] = 46117;
mem_k_index[9872] = 46120;
mem_k_index[9873] = 46122;
mem_k_index[9874] = 46125;
mem_k_index[9875] = 46127;
mem_k_index[9876] = 46130;
mem_k_index[9877] = 46132;
mem_k_index[9878] = 46135;
mem_k_index[9879] = 46137;
mem_k_index[9880] = 46140;
mem_k_index[9881] = 46142;
mem_k_index[9882] = 46145;
mem_k_index[9883] = 46147;
mem_k_index[9884] = 46150;
mem_k_index[9885] = 46152;
mem_k_index[9886] = 46155;
mem_k_index[9887] = 46157;
mem_k_index[9888] = 46160;
mem_k_index[9889] = 46162;
mem_k_index[9890] = 46165;
mem_k_index[9891] = 46167;
mem_k_index[9892] = 46170;
mem_k_index[9893] = 46172;
mem_k_index[9894] = 46175;
mem_k_index[9895] = 46177;
mem_k_index[9896] = 46180;
mem_k_index[9897] = 46182;
mem_k_index[9898] = 46185;
mem_k_index[9899] = 46188;
mem_k_index[9900] = 46190;
mem_k_index[9901] = 46193;
mem_k_index[9902] = 46195;
mem_k_index[9903] = 46198;
mem_k_index[9904] = 46200;
mem_k_index[9905] = 46203;
mem_k_index[9906] = 46205;
mem_k_index[9907] = 46208;
mem_k_index[9908] = 46210;
mem_k_index[9909] = 46213;
mem_k_index[9910] = 46215;
mem_k_index[9911] = 46218;
mem_k_index[9912] = 46220;
mem_k_index[9913] = 46223;
mem_k_index[9914] = 46225;
mem_k_index[9915] = 46228;
mem_k_index[9916] = 46230;
mem_k_index[9917] = 46233;
mem_k_index[9918] = 46235;
mem_k_index[9919] = 46238;
mem_k_index[9920] = 46240;
mem_k_index[9921] = 46243;
mem_k_index[9922] = 46245;
mem_k_index[9923] = 46248;
mem_k_index[9924] = 46250;
mem_k_index[9925] = 46253;
mem_k_index[9926] = 46255;
mem_k_index[9927] = 46258;
mem_k_index[9928] = 46260;
mem_k_index[9929] = 46263;
mem_k_index[9930] = 46265;
mem_k_index[9931] = 46268;
mem_k_index[9932] = 46270;
mem_k_index[9933] = 46273;
mem_k_index[9934] = 46275;
mem_k_index[9935] = 46278;
mem_k_index[9936] = 46280;
mem_k_index[9937] = 46283;
mem_k_index[9938] = 46285;
mem_k_index[9939] = 46288;
mem_k_index[9940] = 46290;
mem_k_index[9941] = 46293;
mem_k_index[9942] = 46296;
mem_k_index[9943] = 46298;
mem_k_index[9944] = 46301;
mem_k_index[9945] = 46303;
mem_k_index[9946] = 46306;
mem_k_index[9947] = 46308;
mem_k_index[9948] = 46311;
mem_k_index[9949] = 46313;
mem_k_index[9950] = 46316;
mem_k_index[9951] = 46318;
mem_k_index[9952] = 46321;
mem_k_index[9953] = 46323;
mem_k_index[9954] = 46326;
mem_k_index[9955] = 46328;
mem_k_index[9956] = 46331;
mem_k_index[9957] = 46333;
mem_k_index[9958] = 46336;
mem_k_index[9959] = 46338;
mem_k_index[9960] = 46341;
mem_k_index[9961] = 46343;
mem_k_index[9962] = 46346;
mem_k_index[9963] = 46348;
mem_k_index[9964] = 46351;
mem_k_index[9965] = 46353;
mem_k_index[9966] = 46356;
mem_k_index[9967] = 46358;
mem_k_index[9968] = 46361;
mem_k_index[9969] = 46363;
mem_k_index[9970] = 46366;
mem_k_index[9971] = 46368;
mem_k_index[9972] = 46371;
mem_k_index[9973] = 46373;
mem_k_index[9974] = 46376;
mem_k_index[9975] = 46378;
mem_k_index[9976] = 46381;
mem_k_index[9977] = 46383;
mem_k_index[9978] = 46386;
mem_k_index[9979] = 46388;
mem_k_index[9980] = 46391;
mem_k_index[9981] = 46393;
mem_k_index[9982] = 46396;
mem_k_index[9983] = 46398;
mem_k_index[9984] = 46720;
mem_k_index[9985] = 46722;
mem_k_index[9986] = 46725;
mem_k_index[9987] = 46727;
mem_k_index[9988] = 46730;
mem_k_index[9989] = 46732;
mem_k_index[9990] = 46735;
mem_k_index[9991] = 46737;
mem_k_index[9992] = 46740;
mem_k_index[9993] = 46742;
mem_k_index[9994] = 46745;
mem_k_index[9995] = 46747;
mem_k_index[9996] = 46750;
mem_k_index[9997] = 46752;
mem_k_index[9998] = 46755;
mem_k_index[9999] = 46757;
mem_k_index[10000] = 46760;
mem_k_index[10001] = 46762;
mem_k_index[10002] = 46765;
mem_k_index[10003] = 46767;
mem_k_index[10004] = 46770;
mem_k_index[10005] = 46772;
mem_k_index[10006] = 46775;
mem_k_index[10007] = 46777;
mem_k_index[10008] = 46780;
mem_k_index[10009] = 46782;
mem_k_index[10010] = 46785;
mem_k_index[10011] = 46787;
mem_k_index[10012] = 46790;
mem_k_index[10013] = 46792;
mem_k_index[10014] = 46795;
mem_k_index[10015] = 46797;
mem_k_index[10016] = 46800;
mem_k_index[10017] = 46802;
mem_k_index[10018] = 46805;
mem_k_index[10019] = 46807;
mem_k_index[10020] = 46810;
mem_k_index[10021] = 46812;
mem_k_index[10022] = 46815;
mem_k_index[10023] = 46817;
mem_k_index[10024] = 46820;
mem_k_index[10025] = 46822;
mem_k_index[10026] = 46825;
mem_k_index[10027] = 46828;
mem_k_index[10028] = 46830;
mem_k_index[10029] = 46833;
mem_k_index[10030] = 46835;
mem_k_index[10031] = 46838;
mem_k_index[10032] = 46840;
mem_k_index[10033] = 46843;
mem_k_index[10034] = 46845;
mem_k_index[10035] = 46848;
mem_k_index[10036] = 46850;
mem_k_index[10037] = 46853;
mem_k_index[10038] = 46855;
mem_k_index[10039] = 46858;
mem_k_index[10040] = 46860;
mem_k_index[10041] = 46863;
mem_k_index[10042] = 46865;
mem_k_index[10043] = 46868;
mem_k_index[10044] = 46870;
mem_k_index[10045] = 46873;
mem_k_index[10046] = 46875;
mem_k_index[10047] = 46878;
mem_k_index[10048] = 46880;
mem_k_index[10049] = 46883;
mem_k_index[10050] = 46885;
mem_k_index[10051] = 46888;
mem_k_index[10052] = 46890;
mem_k_index[10053] = 46893;
mem_k_index[10054] = 46895;
mem_k_index[10055] = 46898;
mem_k_index[10056] = 46900;
mem_k_index[10057] = 46903;
mem_k_index[10058] = 46905;
mem_k_index[10059] = 46908;
mem_k_index[10060] = 46910;
mem_k_index[10061] = 46913;
mem_k_index[10062] = 46915;
mem_k_index[10063] = 46918;
mem_k_index[10064] = 46920;
mem_k_index[10065] = 46923;
mem_k_index[10066] = 46925;
mem_k_index[10067] = 46928;
mem_k_index[10068] = 46930;
mem_k_index[10069] = 46933;
mem_k_index[10070] = 46936;
mem_k_index[10071] = 46938;
mem_k_index[10072] = 46941;
mem_k_index[10073] = 46943;
mem_k_index[10074] = 46946;
mem_k_index[10075] = 46948;
mem_k_index[10076] = 46951;
mem_k_index[10077] = 46953;
mem_k_index[10078] = 46956;
mem_k_index[10079] = 46958;
mem_k_index[10080] = 46961;
mem_k_index[10081] = 46963;
mem_k_index[10082] = 46966;
mem_k_index[10083] = 46968;
mem_k_index[10084] = 46971;
mem_k_index[10085] = 46973;
mem_k_index[10086] = 46976;
mem_k_index[10087] = 46978;
mem_k_index[10088] = 46981;
mem_k_index[10089] = 46983;
mem_k_index[10090] = 46986;
mem_k_index[10091] = 46988;
mem_k_index[10092] = 46991;
mem_k_index[10093] = 46993;
mem_k_index[10094] = 46996;
mem_k_index[10095] = 46998;
mem_k_index[10096] = 47001;
mem_k_index[10097] = 47003;
mem_k_index[10098] = 47006;
mem_k_index[10099] = 47008;
mem_k_index[10100] = 47011;
mem_k_index[10101] = 47013;
mem_k_index[10102] = 47016;
mem_k_index[10103] = 47018;
mem_k_index[10104] = 47021;
mem_k_index[10105] = 47023;
mem_k_index[10106] = 47026;
mem_k_index[10107] = 47028;
mem_k_index[10108] = 47031;
mem_k_index[10109] = 47033;
mem_k_index[10110] = 47036;
mem_k_index[10111] = 47038;
mem_k_index[10112] = 47360;
mem_k_index[10113] = 47362;
mem_k_index[10114] = 47365;
mem_k_index[10115] = 47367;
mem_k_index[10116] = 47370;
mem_k_index[10117] = 47372;
mem_k_index[10118] = 47375;
mem_k_index[10119] = 47377;
mem_k_index[10120] = 47380;
mem_k_index[10121] = 47382;
mem_k_index[10122] = 47385;
mem_k_index[10123] = 47387;
mem_k_index[10124] = 47390;
mem_k_index[10125] = 47392;
mem_k_index[10126] = 47395;
mem_k_index[10127] = 47397;
mem_k_index[10128] = 47400;
mem_k_index[10129] = 47402;
mem_k_index[10130] = 47405;
mem_k_index[10131] = 47407;
mem_k_index[10132] = 47410;
mem_k_index[10133] = 47412;
mem_k_index[10134] = 47415;
mem_k_index[10135] = 47417;
mem_k_index[10136] = 47420;
mem_k_index[10137] = 47422;
mem_k_index[10138] = 47425;
mem_k_index[10139] = 47427;
mem_k_index[10140] = 47430;
mem_k_index[10141] = 47432;
mem_k_index[10142] = 47435;
mem_k_index[10143] = 47437;
mem_k_index[10144] = 47440;
mem_k_index[10145] = 47442;
mem_k_index[10146] = 47445;
mem_k_index[10147] = 47447;
mem_k_index[10148] = 47450;
mem_k_index[10149] = 47452;
mem_k_index[10150] = 47455;
mem_k_index[10151] = 47457;
mem_k_index[10152] = 47460;
mem_k_index[10153] = 47462;
mem_k_index[10154] = 47465;
mem_k_index[10155] = 47468;
mem_k_index[10156] = 47470;
mem_k_index[10157] = 47473;
mem_k_index[10158] = 47475;
mem_k_index[10159] = 47478;
mem_k_index[10160] = 47480;
mem_k_index[10161] = 47483;
mem_k_index[10162] = 47485;
mem_k_index[10163] = 47488;
mem_k_index[10164] = 47490;
mem_k_index[10165] = 47493;
mem_k_index[10166] = 47495;
mem_k_index[10167] = 47498;
mem_k_index[10168] = 47500;
mem_k_index[10169] = 47503;
mem_k_index[10170] = 47505;
mem_k_index[10171] = 47508;
mem_k_index[10172] = 47510;
mem_k_index[10173] = 47513;
mem_k_index[10174] = 47515;
mem_k_index[10175] = 47518;
mem_k_index[10176] = 47520;
mem_k_index[10177] = 47523;
mem_k_index[10178] = 47525;
mem_k_index[10179] = 47528;
mem_k_index[10180] = 47530;
mem_k_index[10181] = 47533;
mem_k_index[10182] = 47535;
mem_k_index[10183] = 47538;
mem_k_index[10184] = 47540;
mem_k_index[10185] = 47543;
mem_k_index[10186] = 47545;
mem_k_index[10187] = 47548;
mem_k_index[10188] = 47550;
mem_k_index[10189] = 47553;
mem_k_index[10190] = 47555;
mem_k_index[10191] = 47558;
mem_k_index[10192] = 47560;
mem_k_index[10193] = 47563;
mem_k_index[10194] = 47565;
mem_k_index[10195] = 47568;
mem_k_index[10196] = 47570;
mem_k_index[10197] = 47573;
mem_k_index[10198] = 47576;
mem_k_index[10199] = 47578;
mem_k_index[10200] = 47581;
mem_k_index[10201] = 47583;
mem_k_index[10202] = 47586;
mem_k_index[10203] = 47588;
mem_k_index[10204] = 47591;
mem_k_index[10205] = 47593;
mem_k_index[10206] = 47596;
mem_k_index[10207] = 47598;
mem_k_index[10208] = 47601;
mem_k_index[10209] = 47603;
mem_k_index[10210] = 47606;
mem_k_index[10211] = 47608;
mem_k_index[10212] = 47611;
mem_k_index[10213] = 47613;
mem_k_index[10214] = 47616;
mem_k_index[10215] = 47618;
mem_k_index[10216] = 47621;
mem_k_index[10217] = 47623;
mem_k_index[10218] = 47626;
mem_k_index[10219] = 47628;
mem_k_index[10220] = 47631;
mem_k_index[10221] = 47633;
mem_k_index[10222] = 47636;
mem_k_index[10223] = 47638;
mem_k_index[10224] = 47641;
mem_k_index[10225] = 47643;
mem_k_index[10226] = 47646;
mem_k_index[10227] = 47648;
mem_k_index[10228] = 47651;
mem_k_index[10229] = 47653;
mem_k_index[10230] = 47656;
mem_k_index[10231] = 47658;
mem_k_index[10232] = 47661;
mem_k_index[10233] = 47663;
mem_k_index[10234] = 47666;
mem_k_index[10235] = 47668;
mem_k_index[10236] = 47671;
mem_k_index[10237] = 47673;
mem_k_index[10238] = 47676;
mem_k_index[10239] = 47678;
mem_k_index[10240] = 48000;
mem_k_index[10241] = 48002;
mem_k_index[10242] = 48005;
mem_k_index[10243] = 48007;
mem_k_index[10244] = 48010;
mem_k_index[10245] = 48012;
mem_k_index[10246] = 48015;
mem_k_index[10247] = 48017;
mem_k_index[10248] = 48020;
mem_k_index[10249] = 48022;
mem_k_index[10250] = 48025;
mem_k_index[10251] = 48027;
mem_k_index[10252] = 48030;
mem_k_index[10253] = 48032;
mem_k_index[10254] = 48035;
mem_k_index[10255] = 48037;
mem_k_index[10256] = 48040;
mem_k_index[10257] = 48042;
mem_k_index[10258] = 48045;
mem_k_index[10259] = 48047;
mem_k_index[10260] = 48050;
mem_k_index[10261] = 48052;
mem_k_index[10262] = 48055;
mem_k_index[10263] = 48057;
mem_k_index[10264] = 48060;
mem_k_index[10265] = 48062;
mem_k_index[10266] = 48065;
mem_k_index[10267] = 48067;
mem_k_index[10268] = 48070;
mem_k_index[10269] = 48072;
mem_k_index[10270] = 48075;
mem_k_index[10271] = 48077;
mem_k_index[10272] = 48080;
mem_k_index[10273] = 48082;
mem_k_index[10274] = 48085;
mem_k_index[10275] = 48087;
mem_k_index[10276] = 48090;
mem_k_index[10277] = 48092;
mem_k_index[10278] = 48095;
mem_k_index[10279] = 48097;
mem_k_index[10280] = 48100;
mem_k_index[10281] = 48102;
mem_k_index[10282] = 48105;
mem_k_index[10283] = 48108;
mem_k_index[10284] = 48110;
mem_k_index[10285] = 48113;
mem_k_index[10286] = 48115;
mem_k_index[10287] = 48118;
mem_k_index[10288] = 48120;
mem_k_index[10289] = 48123;
mem_k_index[10290] = 48125;
mem_k_index[10291] = 48128;
mem_k_index[10292] = 48130;
mem_k_index[10293] = 48133;
mem_k_index[10294] = 48135;
mem_k_index[10295] = 48138;
mem_k_index[10296] = 48140;
mem_k_index[10297] = 48143;
mem_k_index[10298] = 48145;
mem_k_index[10299] = 48148;
mem_k_index[10300] = 48150;
mem_k_index[10301] = 48153;
mem_k_index[10302] = 48155;
mem_k_index[10303] = 48158;
mem_k_index[10304] = 48160;
mem_k_index[10305] = 48163;
mem_k_index[10306] = 48165;
mem_k_index[10307] = 48168;
mem_k_index[10308] = 48170;
mem_k_index[10309] = 48173;
mem_k_index[10310] = 48175;
mem_k_index[10311] = 48178;
mem_k_index[10312] = 48180;
mem_k_index[10313] = 48183;
mem_k_index[10314] = 48185;
mem_k_index[10315] = 48188;
mem_k_index[10316] = 48190;
mem_k_index[10317] = 48193;
mem_k_index[10318] = 48195;
mem_k_index[10319] = 48198;
mem_k_index[10320] = 48200;
mem_k_index[10321] = 48203;
mem_k_index[10322] = 48205;
mem_k_index[10323] = 48208;
mem_k_index[10324] = 48210;
mem_k_index[10325] = 48213;
mem_k_index[10326] = 48216;
mem_k_index[10327] = 48218;
mem_k_index[10328] = 48221;
mem_k_index[10329] = 48223;
mem_k_index[10330] = 48226;
mem_k_index[10331] = 48228;
mem_k_index[10332] = 48231;
mem_k_index[10333] = 48233;
mem_k_index[10334] = 48236;
mem_k_index[10335] = 48238;
mem_k_index[10336] = 48241;
mem_k_index[10337] = 48243;
mem_k_index[10338] = 48246;
mem_k_index[10339] = 48248;
mem_k_index[10340] = 48251;
mem_k_index[10341] = 48253;
mem_k_index[10342] = 48256;
mem_k_index[10343] = 48258;
mem_k_index[10344] = 48261;
mem_k_index[10345] = 48263;
mem_k_index[10346] = 48266;
mem_k_index[10347] = 48268;
mem_k_index[10348] = 48271;
mem_k_index[10349] = 48273;
mem_k_index[10350] = 48276;
mem_k_index[10351] = 48278;
mem_k_index[10352] = 48281;
mem_k_index[10353] = 48283;
mem_k_index[10354] = 48286;
mem_k_index[10355] = 48288;
mem_k_index[10356] = 48291;
mem_k_index[10357] = 48293;
mem_k_index[10358] = 48296;
mem_k_index[10359] = 48298;
mem_k_index[10360] = 48301;
mem_k_index[10361] = 48303;
mem_k_index[10362] = 48306;
mem_k_index[10363] = 48308;
mem_k_index[10364] = 48311;
mem_k_index[10365] = 48313;
mem_k_index[10366] = 48316;
mem_k_index[10367] = 48318;
mem_k_index[10368] = 48640;
mem_k_index[10369] = 48642;
mem_k_index[10370] = 48645;
mem_k_index[10371] = 48647;
mem_k_index[10372] = 48650;
mem_k_index[10373] = 48652;
mem_k_index[10374] = 48655;
mem_k_index[10375] = 48657;
mem_k_index[10376] = 48660;
mem_k_index[10377] = 48662;
mem_k_index[10378] = 48665;
mem_k_index[10379] = 48667;
mem_k_index[10380] = 48670;
mem_k_index[10381] = 48672;
mem_k_index[10382] = 48675;
mem_k_index[10383] = 48677;
mem_k_index[10384] = 48680;
mem_k_index[10385] = 48682;
mem_k_index[10386] = 48685;
mem_k_index[10387] = 48687;
mem_k_index[10388] = 48690;
mem_k_index[10389] = 48692;
mem_k_index[10390] = 48695;
mem_k_index[10391] = 48697;
mem_k_index[10392] = 48700;
mem_k_index[10393] = 48702;
mem_k_index[10394] = 48705;
mem_k_index[10395] = 48707;
mem_k_index[10396] = 48710;
mem_k_index[10397] = 48712;
mem_k_index[10398] = 48715;
mem_k_index[10399] = 48717;
mem_k_index[10400] = 48720;
mem_k_index[10401] = 48722;
mem_k_index[10402] = 48725;
mem_k_index[10403] = 48727;
mem_k_index[10404] = 48730;
mem_k_index[10405] = 48732;
mem_k_index[10406] = 48735;
mem_k_index[10407] = 48737;
mem_k_index[10408] = 48740;
mem_k_index[10409] = 48742;
mem_k_index[10410] = 48745;
mem_k_index[10411] = 48748;
mem_k_index[10412] = 48750;
mem_k_index[10413] = 48753;
mem_k_index[10414] = 48755;
mem_k_index[10415] = 48758;
mem_k_index[10416] = 48760;
mem_k_index[10417] = 48763;
mem_k_index[10418] = 48765;
mem_k_index[10419] = 48768;
mem_k_index[10420] = 48770;
mem_k_index[10421] = 48773;
mem_k_index[10422] = 48775;
mem_k_index[10423] = 48778;
mem_k_index[10424] = 48780;
mem_k_index[10425] = 48783;
mem_k_index[10426] = 48785;
mem_k_index[10427] = 48788;
mem_k_index[10428] = 48790;
mem_k_index[10429] = 48793;
mem_k_index[10430] = 48795;
mem_k_index[10431] = 48798;
mem_k_index[10432] = 48800;
mem_k_index[10433] = 48803;
mem_k_index[10434] = 48805;
mem_k_index[10435] = 48808;
mem_k_index[10436] = 48810;
mem_k_index[10437] = 48813;
mem_k_index[10438] = 48815;
mem_k_index[10439] = 48818;
mem_k_index[10440] = 48820;
mem_k_index[10441] = 48823;
mem_k_index[10442] = 48825;
mem_k_index[10443] = 48828;
mem_k_index[10444] = 48830;
mem_k_index[10445] = 48833;
mem_k_index[10446] = 48835;
mem_k_index[10447] = 48838;
mem_k_index[10448] = 48840;
mem_k_index[10449] = 48843;
mem_k_index[10450] = 48845;
mem_k_index[10451] = 48848;
mem_k_index[10452] = 48850;
mem_k_index[10453] = 48853;
mem_k_index[10454] = 48856;
mem_k_index[10455] = 48858;
mem_k_index[10456] = 48861;
mem_k_index[10457] = 48863;
mem_k_index[10458] = 48866;
mem_k_index[10459] = 48868;
mem_k_index[10460] = 48871;
mem_k_index[10461] = 48873;
mem_k_index[10462] = 48876;
mem_k_index[10463] = 48878;
mem_k_index[10464] = 48881;
mem_k_index[10465] = 48883;
mem_k_index[10466] = 48886;
mem_k_index[10467] = 48888;
mem_k_index[10468] = 48891;
mem_k_index[10469] = 48893;
mem_k_index[10470] = 48896;
mem_k_index[10471] = 48898;
mem_k_index[10472] = 48901;
mem_k_index[10473] = 48903;
mem_k_index[10474] = 48906;
mem_k_index[10475] = 48908;
mem_k_index[10476] = 48911;
mem_k_index[10477] = 48913;
mem_k_index[10478] = 48916;
mem_k_index[10479] = 48918;
mem_k_index[10480] = 48921;
mem_k_index[10481] = 48923;
mem_k_index[10482] = 48926;
mem_k_index[10483] = 48928;
mem_k_index[10484] = 48931;
mem_k_index[10485] = 48933;
mem_k_index[10486] = 48936;
mem_k_index[10487] = 48938;
mem_k_index[10488] = 48941;
mem_k_index[10489] = 48943;
mem_k_index[10490] = 48946;
mem_k_index[10491] = 48948;
mem_k_index[10492] = 48951;
mem_k_index[10493] = 48953;
mem_k_index[10494] = 48956;
mem_k_index[10495] = 48958;
mem_k_index[10496] = 49280;
mem_k_index[10497] = 49282;
mem_k_index[10498] = 49285;
mem_k_index[10499] = 49287;
mem_k_index[10500] = 49290;
mem_k_index[10501] = 49292;
mem_k_index[10502] = 49295;
mem_k_index[10503] = 49297;
mem_k_index[10504] = 49300;
mem_k_index[10505] = 49302;
mem_k_index[10506] = 49305;
mem_k_index[10507] = 49307;
mem_k_index[10508] = 49310;
mem_k_index[10509] = 49312;
mem_k_index[10510] = 49315;
mem_k_index[10511] = 49317;
mem_k_index[10512] = 49320;
mem_k_index[10513] = 49322;
mem_k_index[10514] = 49325;
mem_k_index[10515] = 49327;
mem_k_index[10516] = 49330;
mem_k_index[10517] = 49332;
mem_k_index[10518] = 49335;
mem_k_index[10519] = 49337;
mem_k_index[10520] = 49340;
mem_k_index[10521] = 49342;
mem_k_index[10522] = 49345;
mem_k_index[10523] = 49347;
mem_k_index[10524] = 49350;
mem_k_index[10525] = 49352;
mem_k_index[10526] = 49355;
mem_k_index[10527] = 49357;
mem_k_index[10528] = 49360;
mem_k_index[10529] = 49362;
mem_k_index[10530] = 49365;
mem_k_index[10531] = 49367;
mem_k_index[10532] = 49370;
mem_k_index[10533] = 49372;
mem_k_index[10534] = 49375;
mem_k_index[10535] = 49377;
mem_k_index[10536] = 49380;
mem_k_index[10537] = 49382;
mem_k_index[10538] = 49385;
mem_k_index[10539] = 49388;
mem_k_index[10540] = 49390;
mem_k_index[10541] = 49393;
mem_k_index[10542] = 49395;
mem_k_index[10543] = 49398;
mem_k_index[10544] = 49400;
mem_k_index[10545] = 49403;
mem_k_index[10546] = 49405;
mem_k_index[10547] = 49408;
mem_k_index[10548] = 49410;
mem_k_index[10549] = 49413;
mem_k_index[10550] = 49415;
mem_k_index[10551] = 49418;
mem_k_index[10552] = 49420;
mem_k_index[10553] = 49423;
mem_k_index[10554] = 49425;
mem_k_index[10555] = 49428;
mem_k_index[10556] = 49430;
mem_k_index[10557] = 49433;
mem_k_index[10558] = 49435;
mem_k_index[10559] = 49438;
mem_k_index[10560] = 49440;
mem_k_index[10561] = 49443;
mem_k_index[10562] = 49445;
mem_k_index[10563] = 49448;
mem_k_index[10564] = 49450;
mem_k_index[10565] = 49453;
mem_k_index[10566] = 49455;
mem_k_index[10567] = 49458;
mem_k_index[10568] = 49460;
mem_k_index[10569] = 49463;
mem_k_index[10570] = 49465;
mem_k_index[10571] = 49468;
mem_k_index[10572] = 49470;
mem_k_index[10573] = 49473;
mem_k_index[10574] = 49475;
mem_k_index[10575] = 49478;
mem_k_index[10576] = 49480;
mem_k_index[10577] = 49483;
mem_k_index[10578] = 49485;
mem_k_index[10579] = 49488;
mem_k_index[10580] = 49490;
mem_k_index[10581] = 49493;
mem_k_index[10582] = 49496;
mem_k_index[10583] = 49498;
mem_k_index[10584] = 49501;
mem_k_index[10585] = 49503;
mem_k_index[10586] = 49506;
mem_k_index[10587] = 49508;
mem_k_index[10588] = 49511;
mem_k_index[10589] = 49513;
mem_k_index[10590] = 49516;
mem_k_index[10591] = 49518;
mem_k_index[10592] = 49521;
mem_k_index[10593] = 49523;
mem_k_index[10594] = 49526;
mem_k_index[10595] = 49528;
mem_k_index[10596] = 49531;
mem_k_index[10597] = 49533;
mem_k_index[10598] = 49536;
mem_k_index[10599] = 49538;
mem_k_index[10600] = 49541;
mem_k_index[10601] = 49543;
mem_k_index[10602] = 49546;
mem_k_index[10603] = 49548;
mem_k_index[10604] = 49551;
mem_k_index[10605] = 49553;
mem_k_index[10606] = 49556;
mem_k_index[10607] = 49558;
mem_k_index[10608] = 49561;
mem_k_index[10609] = 49563;
mem_k_index[10610] = 49566;
mem_k_index[10611] = 49568;
mem_k_index[10612] = 49571;
mem_k_index[10613] = 49573;
mem_k_index[10614] = 49576;
mem_k_index[10615] = 49578;
mem_k_index[10616] = 49581;
mem_k_index[10617] = 49583;
mem_k_index[10618] = 49586;
mem_k_index[10619] = 49588;
mem_k_index[10620] = 49591;
mem_k_index[10621] = 49593;
mem_k_index[10622] = 49596;
mem_k_index[10623] = 49598;
mem_k_index[10624] = 49920;
mem_k_index[10625] = 49922;
mem_k_index[10626] = 49925;
mem_k_index[10627] = 49927;
mem_k_index[10628] = 49930;
mem_k_index[10629] = 49932;
mem_k_index[10630] = 49935;
mem_k_index[10631] = 49937;
mem_k_index[10632] = 49940;
mem_k_index[10633] = 49942;
mem_k_index[10634] = 49945;
mem_k_index[10635] = 49947;
mem_k_index[10636] = 49950;
mem_k_index[10637] = 49952;
mem_k_index[10638] = 49955;
mem_k_index[10639] = 49957;
mem_k_index[10640] = 49960;
mem_k_index[10641] = 49962;
mem_k_index[10642] = 49965;
mem_k_index[10643] = 49967;
mem_k_index[10644] = 49970;
mem_k_index[10645] = 49972;
mem_k_index[10646] = 49975;
mem_k_index[10647] = 49977;
mem_k_index[10648] = 49980;
mem_k_index[10649] = 49982;
mem_k_index[10650] = 49985;
mem_k_index[10651] = 49987;
mem_k_index[10652] = 49990;
mem_k_index[10653] = 49992;
mem_k_index[10654] = 49995;
mem_k_index[10655] = 49997;
mem_k_index[10656] = 50000;
mem_k_index[10657] = 50002;
mem_k_index[10658] = 50005;
mem_k_index[10659] = 50007;
mem_k_index[10660] = 50010;
mem_k_index[10661] = 50012;
mem_k_index[10662] = 50015;
mem_k_index[10663] = 50017;
mem_k_index[10664] = 50020;
mem_k_index[10665] = 50022;
mem_k_index[10666] = 50025;
mem_k_index[10667] = 50028;
mem_k_index[10668] = 50030;
mem_k_index[10669] = 50033;
mem_k_index[10670] = 50035;
mem_k_index[10671] = 50038;
mem_k_index[10672] = 50040;
mem_k_index[10673] = 50043;
mem_k_index[10674] = 50045;
mem_k_index[10675] = 50048;
mem_k_index[10676] = 50050;
mem_k_index[10677] = 50053;
mem_k_index[10678] = 50055;
mem_k_index[10679] = 50058;
mem_k_index[10680] = 50060;
mem_k_index[10681] = 50063;
mem_k_index[10682] = 50065;
mem_k_index[10683] = 50068;
mem_k_index[10684] = 50070;
mem_k_index[10685] = 50073;
mem_k_index[10686] = 50075;
mem_k_index[10687] = 50078;
mem_k_index[10688] = 50080;
mem_k_index[10689] = 50083;
mem_k_index[10690] = 50085;
mem_k_index[10691] = 50088;
mem_k_index[10692] = 50090;
mem_k_index[10693] = 50093;
mem_k_index[10694] = 50095;
mem_k_index[10695] = 50098;
mem_k_index[10696] = 50100;
mem_k_index[10697] = 50103;
mem_k_index[10698] = 50105;
mem_k_index[10699] = 50108;
mem_k_index[10700] = 50110;
mem_k_index[10701] = 50113;
mem_k_index[10702] = 50115;
mem_k_index[10703] = 50118;
mem_k_index[10704] = 50120;
mem_k_index[10705] = 50123;
mem_k_index[10706] = 50125;
mem_k_index[10707] = 50128;
mem_k_index[10708] = 50130;
mem_k_index[10709] = 50133;
mem_k_index[10710] = 50136;
mem_k_index[10711] = 50138;
mem_k_index[10712] = 50141;
mem_k_index[10713] = 50143;
mem_k_index[10714] = 50146;
mem_k_index[10715] = 50148;
mem_k_index[10716] = 50151;
mem_k_index[10717] = 50153;
mem_k_index[10718] = 50156;
mem_k_index[10719] = 50158;
mem_k_index[10720] = 50161;
mem_k_index[10721] = 50163;
mem_k_index[10722] = 50166;
mem_k_index[10723] = 50168;
mem_k_index[10724] = 50171;
mem_k_index[10725] = 50173;
mem_k_index[10726] = 50176;
mem_k_index[10727] = 50178;
mem_k_index[10728] = 50181;
mem_k_index[10729] = 50183;
mem_k_index[10730] = 50186;
mem_k_index[10731] = 50188;
mem_k_index[10732] = 50191;
mem_k_index[10733] = 50193;
mem_k_index[10734] = 50196;
mem_k_index[10735] = 50198;
mem_k_index[10736] = 50201;
mem_k_index[10737] = 50203;
mem_k_index[10738] = 50206;
mem_k_index[10739] = 50208;
mem_k_index[10740] = 50211;
mem_k_index[10741] = 50213;
mem_k_index[10742] = 50216;
mem_k_index[10743] = 50218;
mem_k_index[10744] = 50221;
mem_k_index[10745] = 50223;
mem_k_index[10746] = 50226;
mem_k_index[10747] = 50228;
mem_k_index[10748] = 50231;
mem_k_index[10749] = 50233;
mem_k_index[10750] = 50236;
mem_k_index[10751] = 50238;
mem_k_index[10752] = 50560;
mem_k_index[10753] = 50562;
mem_k_index[10754] = 50565;
mem_k_index[10755] = 50567;
mem_k_index[10756] = 50570;
mem_k_index[10757] = 50572;
mem_k_index[10758] = 50575;
mem_k_index[10759] = 50577;
mem_k_index[10760] = 50580;
mem_k_index[10761] = 50582;
mem_k_index[10762] = 50585;
mem_k_index[10763] = 50587;
mem_k_index[10764] = 50590;
mem_k_index[10765] = 50592;
mem_k_index[10766] = 50595;
mem_k_index[10767] = 50597;
mem_k_index[10768] = 50600;
mem_k_index[10769] = 50602;
mem_k_index[10770] = 50605;
mem_k_index[10771] = 50607;
mem_k_index[10772] = 50610;
mem_k_index[10773] = 50612;
mem_k_index[10774] = 50615;
mem_k_index[10775] = 50617;
mem_k_index[10776] = 50620;
mem_k_index[10777] = 50622;
mem_k_index[10778] = 50625;
mem_k_index[10779] = 50627;
mem_k_index[10780] = 50630;
mem_k_index[10781] = 50632;
mem_k_index[10782] = 50635;
mem_k_index[10783] = 50637;
mem_k_index[10784] = 50640;
mem_k_index[10785] = 50642;
mem_k_index[10786] = 50645;
mem_k_index[10787] = 50647;
mem_k_index[10788] = 50650;
mem_k_index[10789] = 50652;
mem_k_index[10790] = 50655;
mem_k_index[10791] = 50657;
mem_k_index[10792] = 50660;
mem_k_index[10793] = 50662;
mem_k_index[10794] = 50665;
mem_k_index[10795] = 50668;
mem_k_index[10796] = 50670;
mem_k_index[10797] = 50673;
mem_k_index[10798] = 50675;
mem_k_index[10799] = 50678;
mem_k_index[10800] = 50680;
mem_k_index[10801] = 50683;
mem_k_index[10802] = 50685;
mem_k_index[10803] = 50688;
mem_k_index[10804] = 50690;
mem_k_index[10805] = 50693;
mem_k_index[10806] = 50695;
mem_k_index[10807] = 50698;
mem_k_index[10808] = 50700;
mem_k_index[10809] = 50703;
mem_k_index[10810] = 50705;
mem_k_index[10811] = 50708;
mem_k_index[10812] = 50710;
mem_k_index[10813] = 50713;
mem_k_index[10814] = 50715;
mem_k_index[10815] = 50718;
mem_k_index[10816] = 50720;
mem_k_index[10817] = 50723;
mem_k_index[10818] = 50725;
mem_k_index[10819] = 50728;
mem_k_index[10820] = 50730;
mem_k_index[10821] = 50733;
mem_k_index[10822] = 50735;
mem_k_index[10823] = 50738;
mem_k_index[10824] = 50740;
mem_k_index[10825] = 50743;
mem_k_index[10826] = 50745;
mem_k_index[10827] = 50748;
mem_k_index[10828] = 50750;
mem_k_index[10829] = 50753;
mem_k_index[10830] = 50755;
mem_k_index[10831] = 50758;
mem_k_index[10832] = 50760;
mem_k_index[10833] = 50763;
mem_k_index[10834] = 50765;
mem_k_index[10835] = 50768;
mem_k_index[10836] = 50770;
mem_k_index[10837] = 50773;
mem_k_index[10838] = 50776;
mem_k_index[10839] = 50778;
mem_k_index[10840] = 50781;
mem_k_index[10841] = 50783;
mem_k_index[10842] = 50786;
mem_k_index[10843] = 50788;
mem_k_index[10844] = 50791;
mem_k_index[10845] = 50793;
mem_k_index[10846] = 50796;
mem_k_index[10847] = 50798;
mem_k_index[10848] = 50801;
mem_k_index[10849] = 50803;
mem_k_index[10850] = 50806;
mem_k_index[10851] = 50808;
mem_k_index[10852] = 50811;
mem_k_index[10853] = 50813;
mem_k_index[10854] = 50816;
mem_k_index[10855] = 50818;
mem_k_index[10856] = 50821;
mem_k_index[10857] = 50823;
mem_k_index[10858] = 50826;
mem_k_index[10859] = 50828;
mem_k_index[10860] = 50831;
mem_k_index[10861] = 50833;
mem_k_index[10862] = 50836;
mem_k_index[10863] = 50838;
mem_k_index[10864] = 50841;
mem_k_index[10865] = 50843;
mem_k_index[10866] = 50846;
mem_k_index[10867] = 50848;
mem_k_index[10868] = 50851;
mem_k_index[10869] = 50853;
mem_k_index[10870] = 50856;
mem_k_index[10871] = 50858;
mem_k_index[10872] = 50861;
mem_k_index[10873] = 50863;
mem_k_index[10874] = 50866;
mem_k_index[10875] = 50868;
mem_k_index[10876] = 50871;
mem_k_index[10877] = 50873;
mem_k_index[10878] = 50876;
mem_k_index[10879] = 50878;
mem_k_index[10880] = 50880;
mem_k_index[10881] = 50882;
mem_k_index[10882] = 50885;
mem_k_index[10883] = 50887;
mem_k_index[10884] = 50890;
mem_k_index[10885] = 50892;
mem_k_index[10886] = 50895;
mem_k_index[10887] = 50897;
mem_k_index[10888] = 50900;
mem_k_index[10889] = 50902;
mem_k_index[10890] = 50905;
mem_k_index[10891] = 50907;
mem_k_index[10892] = 50910;
mem_k_index[10893] = 50912;
mem_k_index[10894] = 50915;
mem_k_index[10895] = 50917;
mem_k_index[10896] = 50920;
mem_k_index[10897] = 50922;
mem_k_index[10898] = 50925;
mem_k_index[10899] = 50927;
mem_k_index[10900] = 50930;
mem_k_index[10901] = 50932;
mem_k_index[10902] = 50935;
mem_k_index[10903] = 50937;
mem_k_index[10904] = 50940;
mem_k_index[10905] = 50942;
mem_k_index[10906] = 50945;
mem_k_index[10907] = 50947;
mem_k_index[10908] = 50950;
mem_k_index[10909] = 50952;
mem_k_index[10910] = 50955;
mem_k_index[10911] = 50957;
mem_k_index[10912] = 50960;
mem_k_index[10913] = 50962;
mem_k_index[10914] = 50965;
mem_k_index[10915] = 50967;
mem_k_index[10916] = 50970;
mem_k_index[10917] = 50972;
mem_k_index[10918] = 50975;
mem_k_index[10919] = 50977;
mem_k_index[10920] = 50980;
mem_k_index[10921] = 50982;
mem_k_index[10922] = 50985;
mem_k_index[10923] = 50988;
mem_k_index[10924] = 50990;
mem_k_index[10925] = 50993;
mem_k_index[10926] = 50995;
mem_k_index[10927] = 50998;
mem_k_index[10928] = 51000;
mem_k_index[10929] = 51003;
mem_k_index[10930] = 51005;
mem_k_index[10931] = 51008;
mem_k_index[10932] = 51010;
mem_k_index[10933] = 51013;
mem_k_index[10934] = 51015;
mem_k_index[10935] = 51018;
mem_k_index[10936] = 51020;
mem_k_index[10937] = 51023;
mem_k_index[10938] = 51025;
mem_k_index[10939] = 51028;
mem_k_index[10940] = 51030;
mem_k_index[10941] = 51033;
mem_k_index[10942] = 51035;
mem_k_index[10943] = 51038;
mem_k_index[10944] = 51040;
mem_k_index[10945] = 51043;
mem_k_index[10946] = 51045;
mem_k_index[10947] = 51048;
mem_k_index[10948] = 51050;
mem_k_index[10949] = 51053;
mem_k_index[10950] = 51055;
mem_k_index[10951] = 51058;
mem_k_index[10952] = 51060;
mem_k_index[10953] = 51063;
mem_k_index[10954] = 51065;
mem_k_index[10955] = 51068;
mem_k_index[10956] = 51070;
mem_k_index[10957] = 51073;
mem_k_index[10958] = 51075;
mem_k_index[10959] = 51078;
mem_k_index[10960] = 51080;
mem_k_index[10961] = 51083;
mem_k_index[10962] = 51085;
mem_k_index[10963] = 51088;
mem_k_index[10964] = 51090;
mem_k_index[10965] = 51093;
mem_k_index[10966] = 51096;
mem_k_index[10967] = 51098;
mem_k_index[10968] = 51101;
mem_k_index[10969] = 51103;
mem_k_index[10970] = 51106;
mem_k_index[10971] = 51108;
mem_k_index[10972] = 51111;
mem_k_index[10973] = 51113;
mem_k_index[10974] = 51116;
mem_k_index[10975] = 51118;
mem_k_index[10976] = 51121;
mem_k_index[10977] = 51123;
mem_k_index[10978] = 51126;
mem_k_index[10979] = 51128;
mem_k_index[10980] = 51131;
mem_k_index[10981] = 51133;
mem_k_index[10982] = 51136;
mem_k_index[10983] = 51138;
mem_k_index[10984] = 51141;
mem_k_index[10985] = 51143;
mem_k_index[10986] = 51146;
mem_k_index[10987] = 51148;
mem_k_index[10988] = 51151;
mem_k_index[10989] = 51153;
mem_k_index[10990] = 51156;
mem_k_index[10991] = 51158;
mem_k_index[10992] = 51161;
mem_k_index[10993] = 51163;
mem_k_index[10994] = 51166;
mem_k_index[10995] = 51168;
mem_k_index[10996] = 51171;
mem_k_index[10997] = 51173;
mem_k_index[10998] = 51176;
mem_k_index[10999] = 51178;
mem_k_index[11000] = 51181;
mem_k_index[11001] = 51183;
mem_k_index[11002] = 51186;
mem_k_index[11003] = 51188;
mem_k_index[11004] = 51191;
mem_k_index[11005] = 51193;
mem_k_index[11006] = 51196;
mem_k_index[11007] = 51198;
mem_k_index[11008] = 51520;
mem_k_index[11009] = 51522;
mem_k_index[11010] = 51525;
mem_k_index[11011] = 51527;
mem_k_index[11012] = 51530;
mem_k_index[11013] = 51532;
mem_k_index[11014] = 51535;
mem_k_index[11015] = 51537;
mem_k_index[11016] = 51540;
mem_k_index[11017] = 51542;
mem_k_index[11018] = 51545;
mem_k_index[11019] = 51547;
mem_k_index[11020] = 51550;
mem_k_index[11021] = 51552;
mem_k_index[11022] = 51555;
mem_k_index[11023] = 51557;
mem_k_index[11024] = 51560;
mem_k_index[11025] = 51562;
mem_k_index[11026] = 51565;
mem_k_index[11027] = 51567;
mem_k_index[11028] = 51570;
mem_k_index[11029] = 51572;
mem_k_index[11030] = 51575;
mem_k_index[11031] = 51577;
mem_k_index[11032] = 51580;
mem_k_index[11033] = 51582;
mem_k_index[11034] = 51585;
mem_k_index[11035] = 51587;
mem_k_index[11036] = 51590;
mem_k_index[11037] = 51592;
mem_k_index[11038] = 51595;
mem_k_index[11039] = 51597;
mem_k_index[11040] = 51600;
mem_k_index[11041] = 51602;
mem_k_index[11042] = 51605;
mem_k_index[11043] = 51607;
mem_k_index[11044] = 51610;
mem_k_index[11045] = 51612;
mem_k_index[11046] = 51615;
mem_k_index[11047] = 51617;
mem_k_index[11048] = 51620;
mem_k_index[11049] = 51622;
mem_k_index[11050] = 51625;
mem_k_index[11051] = 51628;
mem_k_index[11052] = 51630;
mem_k_index[11053] = 51633;
mem_k_index[11054] = 51635;
mem_k_index[11055] = 51638;
mem_k_index[11056] = 51640;
mem_k_index[11057] = 51643;
mem_k_index[11058] = 51645;
mem_k_index[11059] = 51648;
mem_k_index[11060] = 51650;
mem_k_index[11061] = 51653;
mem_k_index[11062] = 51655;
mem_k_index[11063] = 51658;
mem_k_index[11064] = 51660;
mem_k_index[11065] = 51663;
mem_k_index[11066] = 51665;
mem_k_index[11067] = 51668;
mem_k_index[11068] = 51670;
mem_k_index[11069] = 51673;
mem_k_index[11070] = 51675;
mem_k_index[11071] = 51678;
mem_k_index[11072] = 51680;
mem_k_index[11073] = 51683;
mem_k_index[11074] = 51685;
mem_k_index[11075] = 51688;
mem_k_index[11076] = 51690;
mem_k_index[11077] = 51693;
mem_k_index[11078] = 51695;
mem_k_index[11079] = 51698;
mem_k_index[11080] = 51700;
mem_k_index[11081] = 51703;
mem_k_index[11082] = 51705;
mem_k_index[11083] = 51708;
mem_k_index[11084] = 51710;
mem_k_index[11085] = 51713;
mem_k_index[11086] = 51715;
mem_k_index[11087] = 51718;
mem_k_index[11088] = 51720;
mem_k_index[11089] = 51723;
mem_k_index[11090] = 51725;
mem_k_index[11091] = 51728;
mem_k_index[11092] = 51730;
mem_k_index[11093] = 51733;
mem_k_index[11094] = 51736;
mem_k_index[11095] = 51738;
mem_k_index[11096] = 51741;
mem_k_index[11097] = 51743;
mem_k_index[11098] = 51746;
mem_k_index[11099] = 51748;
mem_k_index[11100] = 51751;
mem_k_index[11101] = 51753;
mem_k_index[11102] = 51756;
mem_k_index[11103] = 51758;
mem_k_index[11104] = 51761;
mem_k_index[11105] = 51763;
mem_k_index[11106] = 51766;
mem_k_index[11107] = 51768;
mem_k_index[11108] = 51771;
mem_k_index[11109] = 51773;
mem_k_index[11110] = 51776;
mem_k_index[11111] = 51778;
mem_k_index[11112] = 51781;
mem_k_index[11113] = 51783;
mem_k_index[11114] = 51786;
mem_k_index[11115] = 51788;
mem_k_index[11116] = 51791;
mem_k_index[11117] = 51793;
mem_k_index[11118] = 51796;
mem_k_index[11119] = 51798;
mem_k_index[11120] = 51801;
mem_k_index[11121] = 51803;
mem_k_index[11122] = 51806;
mem_k_index[11123] = 51808;
mem_k_index[11124] = 51811;
mem_k_index[11125] = 51813;
mem_k_index[11126] = 51816;
mem_k_index[11127] = 51818;
mem_k_index[11128] = 51821;
mem_k_index[11129] = 51823;
mem_k_index[11130] = 51826;
mem_k_index[11131] = 51828;
mem_k_index[11132] = 51831;
mem_k_index[11133] = 51833;
mem_k_index[11134] = 51836;
mem_k_index[11135] = 51838;
mem_k_index[11136] = 52160;
mem_k_index[11137] = 52162;
mem_k_index[11138] = 52165;
mem_k_index[11139] = 52167;
mem_k_index[11140] = 52170;
mem_k_index[11141] = 52172;
mem_k_index[11142] = 52175;
mem_k_index[11143] = 52177;
mem_k_index[11144] = 52180;
mem_k_index[11145] = 52182;
mem_k_index[11146] = 52185;
mem_k_index[11147] = 52187;
mem_k_index[11148] = 52190;
mem_k_index[11149] = 52192;
mem_k_index[11150] = 52195;
mem_k_index[11151] = 52197;
mem_k_index[11152] = 52200;
mem_k_index[11153] = 52202;
mem_k_index[11154] = 52205;
mem_k_index[11155] = 52207;
mem_k_index[11156] = 52210;
mem_k_index[11157] = 52212;
mem_k_index[11158] = 52215;
mem_k_index[11159] = 52217;
mem_k_index[11160] = 52220;
mem_k_index[11161] = 52222;
mem_k_index[11162] = 52225;
mem_k_index[11163] = 52227;
mem_k_index[11164] = 52230;
mem_k_index[11165] = 52232;
mem_k_index[11166] = 52235;
mem_k_index[11167] = 52237;
mem_k_index[11168] = 52240;
mem_k_index[11169] = 52242;
mem_k_index[11170] = 52245;
mem_k_index[11171] = 52247;
mem_k_index[11172] = 52250;
mem_k_index[11173] = 52252;
mem_k_index[11174] = 52255;
mem_k_index[11175] = 52257;
mem_k_index[11176] = 52260;
mem_k_index[11177] = 52262;
mem_k_index[11178] = 52265;
mem_k_index[11179] = 52268;
mem_k_index[11180] = 52270;
mem_k_index[11181] = 52273;
mem_k_index[11182] = 52275;
mem_k_index[11183] = 52278;
mem_k_index[11184] = 52280;
mem_k_index[11185] = 52283;
mem_k_index[11186] = 52285;
mem_k_index[11187] = 52288;
mem_k_index[11188] = 52290;
mem_k_index[11189] = 52293;
mem_k_index[11190] = 52295;
mem_k_index[11191] = 52298;
mem_k_index[11192] = 52300;
mem_k_index[11193] = 52303;
mem_k_index[11194] = 52305;
mem_k_index[11195] = 52308;
mem_k_index[11196] = 52310;
mem_k_index[11197] = 52313;
mem_k_index[11198] = 52315;
mem_k_index[11199] = 52318;
mem_k_index[11200] = 52320;
mem_k_index[11201] = 52323;
mem_k_index[11202] = 52325;
mem_k_index[11203] = 52328;
mem_k_index[11204] = 52330;
mem_k_index[11205] = 52333;
mem_k_index[11206] = 52335;
mem_k_index[11207] = 52338;
mem_k_index[11208] = 52340;
mem_k_index[11209] = 52343;
mem_k_index[11210] = 52345;
mem_k_index[11211] = 52348;
mem_k_index[11212] = 52350;
mem_k_index[11213] = 52353;
mem_k_index[11214] = 52355;
mem_k_index[11215] = 52358;
mem_k_index[11216] = 52360;
mem_k_index[11217] = 52363;
mem_k_index[11218] = 52365;
mem_k_index[11219] = 52368;
mem_k_index[11220] = 52370;
mem_k_index[11221] = 52373;
mem_k_index[11222] = 52376;
mem_k_index[11223] = 52378;
mem_k_index[11224] = 52381;
mem_k_index[11225] = 52383;
mem_k_index[11226] = 52386;
mem_k_index[11227] = 52388;
mem_k_index[11228] = 52391;
mem_k_index[11229] = 52393;
mem_k_index[11230] = 52396;
mem_k_index[11231] = 52398;
mem_k_index[11232] = 52401;
mem_k_index[11233] = 52403;
mem_k_index[11234] = 52406;
mem_k_index[11235] = 52408;
mem_k_index[11236] = 52411;
mem_k_index[11237] = 52413;
mem_k_index[11238] = 52416;
mem_k_index[11239] = 52418;
mem_k_index[11240] = 52421;
mem_k_index[11241] = 52423;
mem_k_index[11242] = 52426;
mem_k_index[11243] = 52428;
mem_k_index[11244] = 52431;
mem_k_index[11245] = 52433;
mem_k_index[11246] = 52436;
mem_k_index[11247] = 52438;
mem_k_index[11248] = 52441;
mem_k_index[11249] = 52443;
mem_k_index[11250] = 52446;
mem_k_index[11251] = 52448;
mem_k_index[11252] = 52451;
mem_k_index[11253] = 52453;
mem_k_index[11254] = 52456;
mem_k_index[11255] = 52458;
mem_k_index[11256] = 52461;
mem_k_index[11257] = 52463;
mem_k_index[11258] = 52466;
mem_k_index[11259] = 52468;
mem_k_index[11260] = 52471;
mem_k_index[11261] = 52473;
mem_k_index[11262] = 52476;
mem_k_index[11263] = 52478;
mem_k_index[11264] = 52800;
mem_k_index[11265] = 52802;
mem_k_index[11266] = 52805;
mem_k_index[11267] = 52807;
mem_k_index[11268] = 52810;
mem_k_index[11269] = 52812;
mem_k_index[11270] = 52815;
mem_k_index[11271] = 52817;
mem_k_index[11272] = 52820;
mem_k_index[11273] = 52822;
mem_k_index[11274] = 52825;
mem_k_index[11275] = 52827;
mem_k_index[11276] = 52830;
mem_k_index[11277] = 52832;
mem_k_index[11278] = 52835;
mem_k_index[11279] = 52837;
mem_k_index[11280] = 52840;
mem_k_index[11281] = 52842;
mem_k_index[11282] = 52845;
mem_k_index[11283] = 52847;
mem_k_index[11284] = 52850;
mem_k_index[11285] = 52852;
mem_k_index[11286] = 52855;
mem_k_index[11287] = 52857;
mem_k_index[11288] = 52860;
mem_k_index[11289] = 52862;
mem_k_index[11290] = 52865;
mem_k_index[11291] = 52867;
mem_k_index[11292] = 52870;
mem_k_index[11293] = 52872;
mem_k_index[11294] = 52875;
mem_k_index[11295] = 52877;
mem_k_index[11296] = 52880;
mem_k_index[11297] = 52882;
mem_k_index[11298] = 52885;
mem_k_index[11299] = 52887;
mem_k_index[11300] = 52890;
mem_k_index[11301] = 52892;
mem_k_index[11302] = 52895;
mem_k_index[11303] = 52897;
mem_k_index[11304] = 52900;
mem_k_index[11305] = 52902;
mem_k_index[11306] = 52905;
mem_k_index[11307] = 52908;
mem_k_index[11308] = 52910;
mem_k_index[11309] = 52913;
mem_k_index[11310] = 52915;
mem_k_index[11311] = 52918;
mem_k_index[11312] = 52920;
mem_k_index[11313] = 52923;
mem_k_index[11314] = 52925;
mem_k_index[11315] = 52928;
mem_k_index[11316] = 52930;
mem_k_index[11317] = 52933;
mem_k_index[11318] = 52935;
mem_k_index[11319] = 52938;
mem_k_index[11320] = 52940;
mem_k_index[11321] = 52943;
mem_k_index[11322] = 52945;
mem_k_index[11323] = 52948;
mem_k_index[11324] = 52950;
mem_k_index[11325] = 52953;
mem_k_index[11326] = 52955;
mem_k_index[11327] = 52958;
mem_k_index[11328] = 52960;
mem_k_index[11329] = 52963;
mem_k_index[11330] = 52965;
mem_k_index[11331] = 52968;
mem_k_index[11332] = 52970;
mem_k_index[11333] = 52973;
mem_k_index[11334] = 52975;
mem_k_index[11335] = 52978;
mem_k_index[11336] = 52980;
mem_k_index[11337] = 52983;
mem_k_index[11338] = 52985;
mem_k_index[11339] = 52988;
mem_k_index[11340] = 52990;
mem_k_index[11341] = 52993;
mem_k_index[11342] = 52995;
mem_k_index[11343] = 52998;
mem_k_index[11344] = 53000;
mem_k_index[11345] = 53003;
mem_k_index[11346] = 53005;
mem_k_index[11347] = 53008;
mem_k_index[11348] = 53010;
mem_k_index[11349] = 53013;
mem_k_index[11350] = 53016;
mem_k_index[11351] = 53018;
mem_k_index[11352] = 53021;
mem_k_index[11353] = 53023;
mem_k_index[11354] = 53026;
mem_k_index[11355] = 53028;
mem_k_index[11356] = 53031;
mem_k_index[11357] = 53033;
mem_k_index[11358] = 53036;
mem_k_index[11359] = 53038;
mem_k_index[11360] = 53041;
mem_k_index[11361] = 53043;
mem_k_index[11362] = 53046;
mem_k_index[11363] = 53048;
mem_k_index[11364] = 53051;
mem_k_index[11365] = 53053;
mem_k_index[11366] = 53056;
mem_k_index[11367] = 53058;
mem_k_index[11368] = 53061;
mem_k_index[11369] = 53063;
mem_k_index[11370] = 53066;
mem_k_index[11371] = 53068;
mem_k_index[11372] = 53071;
mem_k_index[11373] = 53073;
mem_k_index[11374] = 53076;
mem_k_index[11375] = 53078;
mem_k_index[11376] = 53081;
mem_k_index[11377] = 53083;
mem_k_index[11378] = 53086;
mem_k_index[11379] = 53088;
mem_k_index[11380] = 53091;
mem_k_index[11381] = 53093;
mem_k_index[11382] = 53096;
mem_k_index[11383] = 53098;
mem_k_index[11384] = 53101;
mem_k_index[11385] = 53103;
mem_k_index[11386] = 53106;
mem_k_index[11387] = 53108;
mem_k_index[11388] = 53111;
mem_k_index[11389] = 53113;
mem_k_index[11390] = 53116;
mem_k_index[11391] = 53118;
mem_k_index[11392] = 53440;
mem_k_index[11393] = 53442;
mem_k_index[11394] = 53445;
mem_k_index[11395] = 53447;
mem_k_index[11396] = 53450;
mem_k_index[11397] = 53452;
mem_k_index[11398] = 53455;
mem_k_index[11399] = 53457;
mem_k_index[11400] = 53460;
mem_k_index[11401] = 53462;
mem_k_index[11402] = 53465;
mem_k_index[11403] = 53467;
mem_k_index[11404] = 53470;
mem_k_index[11405] = 53472;
mem_k_index[11406] = 53475;
mem_k_index[11407] = 53477;
mem_k_index[11408] = 53480;
mem_k_index[11409] = 53482;
mem_k_index[11410] = 53485;
mem_k_index[11411] = 53487;
mem_k_index[11412] = 53490;
mem_k_index[11413] = 53492;
mem_k_index[11414] = 53495;
mem_k_index[11415] = 53497;
mem_k_index[11416] = 53500;
mem_k_index[11417] = 53502;
mem_k_index[11418] = 53505;
mem_k_index[11419] = 53507;
mem_k_index[11420] = 53510;
mem_k_index[11421] = 53512;
mem_k_index[11422] = 53515;
mem_k_index[11423] = 53517;
mem_k_index[11424] = 53520;
mem_k_index[11425] = 53522;
mem_k_index[11426] = 53525;
mem_k_index[11427] = 53527;
mem_k_index[11428] = 53530;
mem_k_index[11429] = 53532;
mem_k_index[11430] = 53535;
mem_k_index[11431] = 53537;
mem_k_index[11432] = 53540;
mem_k_index[11433] = 53542;
mem_k_index[11434] = 53545;
mem_k_index[11435] = 53548;
mem_k_index[11436] = 53550;
mem_k_index[11437] = 53553;
mem_k_index[11438] = 53555;
mem_k_index[11439] = 53558;
mem_k_index[11440] = 53560;
mem_k_index[11441] = 53563;
mem_k_index[11442] = 53565;
mem_k_index[11443] = 53568;
mem_k_index[11444] = 53570;
mem_k_index[11445] = 53573;
mem_k_index[11446] = 53575;
mem_k_index[11447] = 53578;
mem_k_index[11448] = 53580;
mem_k_index[11449] = 53583;
mem_k_index[11450] = 53585;
mem_k_index[11451] = 53588;
mem_k_index[11452] = 53590;
mem_k_index[11453] = 53593;
mem_k_index[11454] = 53595;
mem_k_index[11455] = 53598;
mem_k_index[11456] = 53600;
mem_k_index[11457] = 53603;
mem_k_index[11458] = 53605;
mem_k_index[11459] = 53608;
mem_k_index[11460] = 53610;
mem_k_index[11461] = 53613;
mem_k_index[11462] = 53615;
mem_k_index[11463] = 53618;
mem_k_index[11464] = 53620;
mem_k_index[11465] = 53623;
mem_k_index[11466] = 53625;
mem_k_index[11467] = 53628;
mem_k_index[11468] = 53630;
mem_k_index[11469] = 53633;
mem_k_index[11470] = 53635;
mem_k_index[11471] = 53638;
mem_k_index[11472] = 53640;
mem_k_index[11473] = 53643;
mem_k_index[11474] = 53645;
mem_k_index[11475] = 53648;
mem_k_index[11476] = 53650;
mem_k_index[11477] = 53653;
mem_k_index[11478] = 53656;
mem_k_index[11479] = 53658;
mem_k_index[11480] = 53661;
mem_k_index[11481] = 53663;
mem_k_index[11482] = 53666;
mem_k_index[11483] = 53668;
mem_k_index[11484] = 53671;
mem_k_index[11485] = 53673;
mem_k_index[11486] = 53676;
mem_k_index[11487] = 53678;
mem_k_index[11488] = 53681;
mem_k_index[11489] = 53683;
mem_k_index[11490] = 53686;
mem_k_index[11491] = 53688;
mem_k_index[11492] = 53691;
mem_k_index[11493] = 53693;
mem_k_index[11494] = 53696;
mem_k_index[11495] = 53698;
mem_k_index[11496] = 53701;
mem_k_index[11497] = 53703;
mem_k_index[11498] = 53706;
mem_k_index[11499] = 53708;
mem_k_index[11500] = 53711;
mem_k_index[11501] = 53713;
mem_k_index[11502] = 53716;
mem_k_index[11503] = 53718;
mem_k_index[11504] = 53721;
mem_k_index[11505] = 53723;
mem_k_index[11506] = 53726;
mem_k_index[11507] = 53728;
mem_k_index[11508] = 53731;
mem_k_index[11509] = 53733;
mem_k_index[11510] = 53736;
mem_k_index[11511] = 53738;
mem_k_index[11512] = 53741;
mem_k_index[11513] = 53743;
mem_k_index[11514] = 53746;
mem_k_index[11515] = 53748;
mem_k_index[11516] = 53751;
mem_k_index[11517] = 53753;
mem_k_index[11518] = 53756;
mem_k_index[11519] = 53758;
mem_k_index[11520] = 54080;
mem_k_index[11521] = 54082;
mem_k_index[11522] = 54085;
mem_k_index[11523] = 54087;
mem_k_index[11524] = 54090;
mem_k_index[11525] = 54092;
mem_k_index[11526] = 54095;
mem_k_index[11527] = 54097;
mem_k_index[11528] = 54100;
mem_k_index[11529] = 54102;
mem_k_index[11530] = 54105;
mem_k_index[11531] = 54107;
mem_k_index[11532] = 54110;
mem_k_index[11533] = 54112;
mem_k_index[11534] = 54115;
mem_k_index[11535] = 54117;
mem_k_index[11536] = 54120;
mem_k_index[11537] = 54122;
mem_k_index[11538] = 54125;
mem_k_index[11539] = 54127;
mem_k_index[11540] = 54130;
mem_k_index[11541] = 54132;
mem_k_index[11542] = 54135;
mem_k_index[11543] = 54137;
mem_k_index[11544] = 54140;
mem_k_index[11545] = 54142;
mem_k_index[11546] = 54145;
mem_k_index[11547] = 54147;
mem_k_index[11548] = 54150;
mem_k_index[11549] = 54152;
mem_k_index[11550] = 54155;
mem_k_index[11551] = 54157;
mem_k_index[11552] = 54160;
mem_k_index[11553] = 54162;
mem_k_index[11554] = 54165;
mem_k_index[11555] = 54167;
mem_k_index[11556] = 54170;
mem_k_index[11557] = 54172;
mem_k_index[11558] = 54175;
mem_k_index[11559] = 54177;
mem_k_index[11560] = 54180;
mem_k_index[11561] = 54182;
mem_k_index[11562] = 54185;
mem_k_index[11563] = 54188;
mem_k_index[11564] = 54190;
mem_k_index[11565] = 54193;
mem_k_index[11566] = 54195;
mem_k_index[11567] = 54198;
mem_k_index[11568] = 54200;
mem_k_index[11569] = 54203;
mem_k_index[11570] = 54205;
mem_k_index[11571] = 54208;
mem_k_index[11572] = 54210;
mem_k_index[11573] = 54213;
mem_k_index[11574] = 54215;
mem_k_index[11575] = 54218;
mem_k_index[11576] = 54220;
mem_k_index[11577] = 54223;
mem_k_index[11578] = 54225;
mem_k_index[11579] = 54228;
mem_k_index[11580] = 54230;
mem_k_index[11581] = 54233;
mem_k_index[11582] = 54235;
mem_k_index[11583] = 54238;
mem_k_index[11584] = 54240;
mem_k_index[11585] = 54243;
mem_k_index[11586] = 54245;
mem_k_index[11587] = 54248;
mem_k_index[11588] = 54250;
mem_k_index[11589] = 54253;
mem_k_index[11590] = 54255;
mem_k_index[11591] = 54258;
mem_k_index[11592] = 54260;
mem_k_index[11593] = 54263;
mem_k_index[11594] = 54265;
mem_k_index[11595] = 54268;
mem_k_index[11596] = 54270;
mem_k_index[11597] = 54273;
mem_k_index[11598] = 54275;
mem_k_index[11599] = 54278;
mem_k_index[11600] = 54280;
mem_k_index[11601] = 54283;
mem_k_index[11602] = 54285;
mem_k_index[11603] = 54288;
mem_k_index[11604] = 54290;
mem_k_index[11605] = 54293;
mem_k_index[11606] = 54296;
mem_k_index[11607] = 54298;
mem_k_index[11608] = 54301;
mem_k_index[11609] = 54303;
mem_k_index[11610] = 54306;
mem_k_index[11611] = 54308;
mem_k_index[11612] = 54311;
mem_k_index[11613] = 54313;
mem_k_index[11614] = 54316;
mem_k_index[11615] = 54318;
mem_k_index[11616] = 54321;
mem_k_index[11617] = 54323;
mem_k_index[11618] = 54326;
mem_k_index[11619] = 54328;
mem_k_index[11620] = 54331;
mem_k_index[11621] = 54333;
mem_k_index[11622] = 54336;
mem_k_index[11623] = 54338;
mem_k_index[11624] = 54341;
mem_k_index[11625] = 54343;
mem_k_index[11626] = 54346;
mem_k_index[11627] = 54348;
mem_k_index[11628] = 54351;
mem_k_index[11629] = 54353;
mem_k_index[11630] = 54356;
mem_k_index[11631] = 54358;
mem_k_index[11632] = 54361;
mem_k_index[11633] = 54363;
mem_k_index[11634] = 54366;
mem_k_index[11635] = 54368;
mem_k_index[11636] = 54371;
mem_k_index[11637] = 54373;
mem_k_index[11638] = 54376;
mem_k_index[11639] = 54378;
mem_k_index[11640] = 54381;
mem_k_index[11641] = 54383;
mem_k_index[11642] = 54386;
mem_k_index[11643] = 54388;
mem_k_index[11644] = 54391;
mem_k_index[11645] = 54393;
mem_k_index[11646] = 54396;
mem_k_index[11647] = 54398;
mem_k_index[11648] = 54720;
mem_k_index[11649] = 54722;
mem_k_index[11650] = 54725;
mem_k_index[11651] = 54727;
mem_k_index[11652] = 54730;
mem_k_index[11653] = 54732;
mem_k_index[11654] = 54735;
mem_k_index[11655] = 54737;
mem_k_index[11656] = 54740;
mem_k_index[11657] = 54742;
mem_k_index[11658] = 54745;
mem_k_index[11659] = 54747;
mem_k_index[11660] = 54750;
mem_k_index[11661] = 54752;
mem_k_index[11662] = 54755;
mem_k_index[11663] = 54757;
mem_k_index[11664] = 54760;
mem_k_index[11665] = 54762;
mem_k_index[11666] = 54765;
mem_k_index[11667] = 54767;
mem_k_index[11668] = 54770;
mem_k_index[11669] = 54772;
mem_k_index[11670] = 54775;
mem_k_index[11671] = 54777;
mem_k_index[11672] = 54780;
mem_k_index[11673] = 54782;
mem_k_index[11674] = 54785;
mem_k_index[11675] = 54787;
mem_k_index[11676] = 54790;
mem_k_index[11677] = 54792;
mem_k_index[11678] = 54795;
mem_k_index[11679] = 54797;
mem_k_index[11680] = 54800;
mem_k_index[11681] = 54802;
mem_k_index[11682] = 54805;
mem_k_index[11683] = 54807;
mem_k_index[11684] = 54810;
mem_k_index[11685] = 54812;
mem_k_index[11686] = 54815;
mem_k_index[11687] = 54817;
mem_k_index[11688] = 54820;
mem_k_index[11689] = 54822;
mem_k_index[11690] = 54825;
mem_k_index[11691] = 54828;
mem_k_index[11692] = 54830;
mem_k_index[11693] = 54833;
mem_k_index[11694] = 54835;
mem_k_index[11695] = 54838;
mem_k_index[11696] = 54840;
mem_k_index[11697] = 54843;
mem_k_index[11698] = 54845;
mem_k_index[11699] = 54848;
mem_k_index[11700] = 54850;
mem_k_index[11701] = 54853;
mem_k_index[11702] = 54855;
mem_k_index[11703] = 54858;
mem_k_index[11704] = 54860;
mem_k_index[11705] = 54863;
mem_k_index[11706] = 54865;
mem_k_index[11707] = 54868;
mem_k_index[11708] = 54870;
mem_k_index[11709] = 54873;
mem_k_index[11710] = 54875;
mem_k_index[11711] = 54878;
mem_k_index[11712] = 54880;
mem_k_index[11713] = 54883;
mem_k_index[11714] = 54885;
mem_k_index[11715] = 54888;
mem_k_index[11716] = 54890;
mem_k_index[11717] = 54893;
mem_k_index[11718] = 54895;
mem_k_index[11719] = 54898;
mem_k_index[11720] = 54900;
mem_k_index[11721] = 54903;
mem_k_index[11722] = 54905;
mem_k_index[11723] = 54908;
mem_k_index[11724] = 54910;
mem_k_index[11725] = 54913;
mem_k_index[11726] = 54915;
mem_k_index[11727] = 54918;
mem_k_index[11728] = 54920;
mem_k_index[11729] = 54923;
mem_k_index[11730] = 54925;
mem_k_index[11731] = 54928;
mem_k_index[11732] = 54930;
mem_k_index[11733] = 54933;
mem_k_index[11734] = 54936;
mem_k_index[11735] = 54938;
mem_k_index[11736] = 54941;
mem_k_index[11737] = 54943;
mem_k_index[11738] = 54946;
mem_k_index[11739] = 54948;
mem_k_index[11740] = 54951;
mem_k_index[11741] = 54953;
mem_k_index[11742] = 54956;
mem_k_index[11743] = 54958;
mem_k_index[11744] = 54961;
mem_k_index[11745] = 54963;
mem_k_index[11746] = 54966;
mem_k_index[11747] = 54968;
mem_k_index[11748] = 54971;
mem_k_index[11749] = 54973;
mem_k_index[11750] = 54976;
mem_k_index[11751] = 54978;
mem_k_index[11752] = 54981;
mem_k_index[11753] = 54983;
mem_k_index[11754] = 54986;
mem_k_index[11755] = 54988;
mem_k_index[11756] = 54991;
mem_k_index[11757] = 54993;
mem_k_index[11758] = 54996;
mem_k_index[11759] = 54998;
mem_k_index[11760] = 55001;
mem_k_index[11761] = 55003;
mem_k_index[11762] = 55006;
mem_k_index[11763] = 55008;
mem_k_index[11764] = 55011;
mem_k_index[11765] = 55013;
mem_k_index[11766] = 55016;
mem_k_index[11767] = 55018;
mem_k_index[11768] = 55021;
mem_k_index[11769] = 55023;
mem_k_index[11770] = 55026;
mem_k_index[11771] = 55028;
mem_k_index[11772] = 55031;
mem_k_index[11773] = 55033;
mem_k_index[11774] = 55036;
mem_k_index[11775] = 55038;
mem_k_index[11776] = 55360;
mem_k_index[11777] = 55362;
mem_k_index[11778] = 55365;
mem_k_index[11779] = 55367;
mem_k_index[11780] = 55370;
mem_k_index[11781] = 55372;
mem_k_index[11782] = 55375;
mem_k_index[11783] = 55377;
mem_k_index[11784] = 55380;
mem_k_index[11785] = 55382;
mem_k_index[11786] = 55385;
mem_k_index[11787] = 55387;
mem_k_index[11788] = 55390;
mem_k_index[11789] = 55392;
mem_k_index[11790] = 55395;
mem_k_index[11791] = 55397;
mem_k_index[11792] = 55400;
mem_k_index[11793] = 55402;
mem_k_index[11794] = 55405;
mem_k_index[11795] = 55407;
mem_k_index[11796] = 55410;
mem_k_index[11797] = 55412;
mem_k_index[11798] = 55415;
mem_k_index[11799] = 55417;
mem_k_index[11800] = 55420;
mem_k_index[11801] = 55422;
mem_k_index[11802] = 55425;
mem_k_index[11803] = 55427;
mem_k_index[11804] = 55430;
mem_k_index[11805] = 55432;
mem_k_index[11806] = 55435;
mem_k_index[11807] = 55437;
mem_k_index[11808] = 55440;
mem_k_index[11809] = 55442;
mem_k_index[11810] = 55445;
mem_k_index[11811] = 55447;
mem_k_index[11812] = 55450;
mem_k_index[11813] = 55452;
mem_k_index[11814] = 55455;
mem_k_index[11815] = 55457;
mem_k_index[11816] = 55460;
mem_k_index[11817] = 55462;
mem_k_index[11818] = 55465;
mem_k_index[11819] = 55468;
mem_k_index[11820] = 55470;
mem_k_index[11821] = 55473;
mem_k_index[11822] = 55475;
mem_k_index[11823] = 55478;
mem_k_index[11824] = 55480;
mem_k_index[11825] = 55483;
mem_k_index[11826] = 55485;
mem_k_index[11827] = 55488;
mem_k_index[11828] = 55490;
mem_k_index[11829] = 55493;
mem_k_index[11830] = 55495;
mem_k_index[11831] = 55498;
mem_k_index[11832] = 55500;
mem_k_index[11833] = 55503;
mem_k_index[11834] = 55505;
mem_k_index[11835] = 55508;
mem_k_index[11836] = 55510;
mem_k_index[11837] = 55513;
mem_k_index[11838] = 55515;
mem_k_index[11839] = 55518;
mem_k_index[11840] = 55520;
mem_k_index[11841] = 55523;
mem_k_index[11842] = 55525;
mem_k_index[11843] = 55528;
mem_k_index[11844] = 55530;
mem_k_index[11845] = 55533;
mem_k_index[11846] = 55535;
mem_k_index[11847] = 55538;
mem_k_index[11848] = 55540;
mem_k_index[11849] = 55543;
mem_k_index[11850] = 55545;
mem_k_index[11851] = 55548;
mem_k_index[11852] = 55550;
mem_k_index[11853] = 55553;
mem_k_index[11854] = 55555;
mem_k_index[11855] = 55558;
mem_k_index[11856] = 55560;
mem_k_index[11857] = 55563;
mem_k_index[11858] = 55565;
mem_k_index[11859] = 55568;
mem_k_index[11860] = 55570;
mem_k_index[11861] = 55573;
mem_k_index[11862] = 55576;
mem_k_index[11863] = 55578;
mem_k_index[11864] = 55581;
mem_k_index[11865] = 55583;
mem_k_index[11866] = 55586;
mem_k_index[11867] = 55588;
mem_k_index[11868] = 55591;
mem_k_index[11869] = 55593;
mem_k_index[11870] = 55596;
mem_k_index[11871] = 55598;
mem_k_index[11872] = 55601;
mem_k_index[11873] = 55603;
mem_k_index[11874] = 55606;
mem_k_index[11875] = 55608;
mem_k_index[11876] = 55611;
mem_k_index[11877] = 55613;
mem_k_index[11878] = 55616;
mem_k_index[11879] = 55618;
mem_k_index[11880] = 55621;
mem_k_index[11881] = 55623;
mem_k_index[11882] = 55626;
mem_k_index[11883] = 55628;
mem_k_index[11884] = 55631;
mem_k_index[11885] = 55633;
mem_k_index[11886] = 55636;
mem_k_index[11887] = 55638;
mem_k_index[11888] = 55641;
mem_k_index[11889] = 55643;
mem_k_index[11890] = 55646;
mem_k_index[11891] = 55648;
mem_k_index[11892] = 55651;
mem_k_index[11893] = 55653;
mem_k_index[11894] = 55656;
mem_k_index[11895] = 55658;
mem_k_index[11896] = 55661;
mem_k_index[11897] = 55663;
mem_k_index[11898] = 55666;
mem_k_index[11899] = 55668;
mem_k_index[11900] = 55671;
mem_k_index[11901] = 55673;
mem_k_index[11902] = 55676;
mem_k_index[11903] = 55678;
mem_k_index[11904] = 56000;
mem_k_index[11905] = 56002;
mem_k_index[11906] = 56005;
mem_k_index[11907] = 56007;
mem_k_index[11908] = 56010;
mem_k_index[11909] = 56012;
mem_k_index[11910] = 56015;
mem_k_index[11911] = 56017;
mem_k_index[11912] = 56020;
mem_k_index[11913] = 56022;
mem_k_index[11914] = 56025;
mem_k_index[11915] = 56027;
mem_k_index[11916] = 56030;
mem_k_index[11917] = 56032;
mem_k_index[11918] = 56035;
mem_k_index[11919] = 56037;
mem_k_index[11920] = 56040;
mem_k_index[11921] = 56042;
mem_k_index[11922] = 56045;
mem_k_index[11923] = 56047;
mem_k_index[11924] = 56050;
mem_k_index[11925] = 56052;
mem_k_index[11926] = 56055;
mem_k_index[11927] = 56057;
mem_k_index[11928] = 56060;
mem_k_index[11929] = 56062;
mem_k_index[11930] = 56065;
mem_k_index[11931] = 56067;
mem_k_index[11932] = 56070;
mem_k_index[11933] = 56072;
mem_k_index[11934] = 56075;
mem_k_index[11935] = 56077;
mem_k_index[11936] = 56080;
mem_k_index[11937] = 56082;
mem_k_index[11938] = 56085;
mem_k_index[11939] = 56087;
mem_k_index[11940] = 56090;
mem_k_index[11941] = 56092;
mem_k_index[11942] = 56095;
mem_k_index[11943] = 56097;
mem_k_index[11944] = 56100;
mem_k_index[11945] = 56102;
mem_k_index[11946] = 56105;
mem_k_index[11947] = 56108;
mem_k_index[11948] = 56110;
mem_k_index[11949] = 56113;
mem_k_index[11950] = 56115;
mem_k_index[11951] = 56118;
mem_k_index[11952] = 56120;
mem_k_index[11953] = 56123;
mem_k_index[11954] = 56125;
mem_k_index[11955] = 56128;
mem_k_index[11956] = 56130;
mem_k_index[11957] = 56133;
mem_k_index[11958] = 56135;
mem_k_index[11959] = 56138;
mem_k_index[11960] = 56140;
mem_k_index[11961] = 56143;
mem_k_index[11962] = 56145;
mem_k_index[11963] = 56148;
mem_k_index[11964] = 56150;
mem_k_index[11965] = 56153;
mem_k_index[11966] = 56155;
mem_k_index[11967] = 56158;
mem_k_index[11968] = 56160;
mem_k_index[11969] = 56163;
mem_k_index[11970] = 56165;
mem_k_index[11971] = 56168;
mem_k_index[11972] = 56170;
mem_k_index[11973] = 56173;
mem_k_index[11974] = 56175;
mem_k_index[11975] = 56178;
mem_k_index[11976] = 56180;
mem_k_index[11977] = 56183;
mem_k_index[11978] = 56185;
mem_k_index[11979] = 56188;
mem_k_index[11980] = 56190;
mem_k_index[11981] = 56193;
mem_k_index[11982] = 56195;
mem_k_index[11983] = 56198;
mem_k_index[11984] = 56200;
mem_k_index[11985] = 56203;
mem_k_index[11986] = 56205;
mem_k_index[11987] = 56208;
mem_k_index[11988] = 56210;
mem_k_index[11989] = 56213;
mem_k_index[11990] = 56216;
mem_k_index[11991] = 56218;
mem_k_index[11992] = 56221;
mem_k_index[11993] = 56223;
mem_k_index[11994] = 56226;
mem_k_index[11995] = 56228;
mem_k_index[11996] = 56231;
mem_k_index[11997] = 56233;
mem_k_index[11998] = 56236;
mem_k_index[11999] = 56238;
mem_k_index[12000] = 56241;
mem_k_index[12001] = 56243;
mem_k_index[12002] = 56246;
mem_k_index[12003] = 56248;
mem_k_index[12004] = 56251;
mem_k_index[12005] = 56253;
mem_k_index[12006] = 56256;
mem_k_index[12007] = 56258;
mem_k_index[12008] = 56261;
mem_k_index[12009] = 56263;
mem_k_index[12010] = 56266;
mem_k_index[12011] = 56268;
mem_k_index[12012] = 56271;
mem_k_index[12013] = 56273;
mem_k_index[12014] = 56276;
mem_k_index[12015] = 56278;
mem_k_index[12016] = 56281;
mem_k_index[12017] = 56283;
mem_k_index[12018] = 56286;
mem_k_index[12019] = 56288;
mem_k_index[12020] = 56291;
mem_k_index[12021] = 56293;
mem_k_index[12022] = 56296;
mem_k_index[12023] = 56298;
mem_k_index[12024] = 56301;
mem_k_index[12025] = 56303;
mem_k_index[12026] = 56306;
mem_k_index[12027] = 56308;
mem_k_index[12028] = 56311;
mem_k_index[12029] = 56313;
mem_k_index[12030] = 56316;
mem_k_index[12031] = 56318;
mem_k_index[12032] = 56320;
mem_k_index[12033] = 56322;
mem_k_index[12034] = 56325;
mem_k_index[12035] = 56327;
mem_k_index[12036] = 56330;
mem_k_index[12037] = 56332;
mem_k_index[12038] = 56335;
mem_k_index[12039] = 56337;
mem_k_index[12040] = 56340;
mem_k_index[12041] = 56342;
mem_k_index[12042] = 56345;
mem_k_index[12043] = 56347;
mem_k_index[12044] = 56350;
mem_k_index[12045] = 56352;
mem_k_index[12046] = 56355;
mem_k_index[12047] = 56357;
mem_k_index[12048] = 56360;
mem_k_index[12049] = 56362;
mem_k_index[12050] = 56365;
mem_k_index[12051] = 56367;
mem_k_index[12052] = 56370;
mem_k_index[12053] = 56372;
mem_k_index[12054] = 56375;
mem_k_index[12055] = 56377;
mem_k_index[12056] = 56380;
mem_k_index[12057] = 56382;
mem_k_index[12058] = 56385;
mem_k_index[12059] = 56387;
mem_k_index[12060] = 56390;
mem_k_index[12061] = 56392;
mem_k_index[12062] = 56395;
mem_k_index[12063] = 56397;
mem_k_index[12064] = 56400;
mem_k_index[12065] = 56402;
mem_k_index[12066] = 56405;
mem_k_index[12067] = 56407;
mem_k_index[12068] = 56410;
mem_k_index[12069] = 56412;
mem_k_index[12070] = 56415;
mem_k_index[12071] = 56417;
mem_k_index[12072] = 56420;
mem_k_index[12073] = 56422;
mem_k_index[12074] = 56425;
mem_k_index[12075] = 56428;
mem_k_index[12076] = 56430;
mem_k_index[12077] = 56433;
mem_k_index[12078] = 56435;
mem_k_index[12079] = 56438;
mem_k_index[12080] = 56440;
mem_k_index[12081] = 56443;
mem_k_index[12082] = 56445;
mem_k_index[12083] = 56448;
mem_k_index[12084] = 56450;
mem_k_index[12085] = 56453;
mem_k_index[12086] = 56455;
mem_k_index[12087] = 56458;
mem_k_index[12088] = 56460;
mem_k_index[12089] = 56463;
mem_k_index[12090] = 56465;
mem_k_index[12091] = 56468;
mem_k_index[12092] = 56470;
mem_k_index[12093] = 56473;
mem_k_index[12094] = 56475;
mem_k_index[12095] = 56478;
mem_k_index[12096] = 56480;
mem_k_index[12097] = 56483;
mem_k_index[12098] = 56485;
mem_k_index[12099] = 56488;
mem_k_index[12100] = 56490;
mem_k_index[12101] = 56493;
mem_k_index[12102] = 56495;
mem_k_index[12103] = 56498;
mem_k_index[12104] = 56500;
mem_k_index[12105] = 56503;
mem_k_index[12106] = 56505;
mem_k_index[12107] = 56508;
mem_k_index[12108] = 56510;
mem_k_index[12109] = 56513;
mem_k_index[12110] = 56515;
mem_k_index[12111] = 56518;
mem_k_index[12112] = 56520;
mem_k_index[12113] = 56523;
mem_k_index[12114] = 56525;
mem_k_index[12115] = 56528;
mem_k_index[12116] = 56530;
mem_k_index[12117] = 56533;
mem_k_index[12118] = 56536;
mem_k_index[12119] = 56538;
mem_k_index[12120] = 56541;
mem_k_index[12121] = 56543;
mem_k_index[12122] = 56546;
mem_k_index[12123] = 56548;
mem_k_index[12124] = 56551;
mem_k_index[12125] = 56553;
mem_k_index[12126] = 56556;
mem_k_index[12127] = 56558;
mem_k_index[12128] = 56561;
mem_k_index[12129] = 56563;
mem_k_index[12130] = 56566;
mem_k_index[12131] = 56568;
mem_k_index[12132] = 56571;
mem_k_index[12133] = 56573;
mem_k_index[12134] = 56576;
mem_k_index[12135] = 56578;
mem_k_index[12136] = 56581;
mem_k_index[12137] = 56583;
mem_k_index[12138] = 56586;
mem_k_index[12139] = 56588;
mem_k_index[12140] = 56591;
mem_k_index[12141] = 56593;
mem_k_index[12142] = 56596;
mem_k_index[12143] = 56598;
mem_k_index[12144] = 56601;
mem_k_index[12145] = 56603;
mem_k_index[12146] = 56606;
mem_k_index[12147] = 56608;
mem_k_index[12148] = 56611;
mem_k_index[12149] = 56613;
mem_k_index[12150] = 56616;
mem_k_index[12151] = 56618;
mem_k_index[12152] = 56621;
mem_k_index[12153] = 56623;
mem_k_index[12154] = 56626;
mem_k_index[12155] = 56628;
mem_k_index[12156] = 56631;
mem_k_index[12157] = 56633;
mem_k_index[12158] = 56636;
mem_k_index[12159] = 56638;
mem_k_index[12160] = 56960;
mem_k_index[12161] = 56962;
mem_k_index[12162] = 56965;
mem_k_index[12163] = 56967;
mem_k_index[12164] = 56970;
mem_k_index[12165] = 56972;
mem_k_index[12166] = 56975;
mem_k_index[12167] = 56977;
mem_k_index[12168] = 56980;
mem_k_index[12169] = 56982;
mem_k_index[12170] = 56985;
mem_k_index[12171] = 56987;
mem_k_index[12172] = 56990;
mem_k_index[12173] = 56992;
mem_k_index[12174] = 56995;
mem_k_index[12175] = 56997;
mem_k_index[12176] = 57000;
mem_k_index[12177] = 57002;
mem_k_index[12178] = 57005;
mem_k_index[12179] = 57007;
mem_k_index[12180] = 57010;
mem_k_index[12181] = 57012;
mem_k_index[12182] = 57015;
mem_k_index[12183] = 57017;
mem_k_index[12184] = 57020;
mem_k_index[12185] = 57022;
mem_k_index[12186] = 57025;
mem_k_index[12187] = 57027;
mem_k_index[12188] = 57030;
mem_k_index[12189] = 57032;
mem_k_index[12190] = 57035;
mem_k_index[12191] = 57037;
mem_k_index[12192] = 57040;
mem_k_index[12193] = 57042;
mem_k_index[12194] = 57045;
mem_k_index[12195] = 57047;
mem_k_index[12196] = 57050;
mem_k_index[12197] = 57052;
mem_k_index[12198] = 57055;
mem_k_index[12199] = 57057;
mem_k_index[12200] = 57060;
mem_k_index[12201] = 57062;
mem_k_index[12202] = 57065;
mem_k_index[12203] = 57068;
mem_k_index[12204] = 57070;
mem_k_index[12205] = 57073;
mem_k_index[12206] = 57075;
mem_k_index[12207] = 57078;
mem_k_index[12208] = 57080;
mem_k_index[12209] = 57083;
mem_k_index[12210] = 57085;
mem_k_index[12211] = 57088;
mem_k_index[12212] = 57090;
mem_k_index[12213] = 57093;
mem_k_index[12214] = 57095;
mem_k_index[12215] = 57098;
mem_k_index[12216] = 57100;
mem_k_index[12217] = 57103;
mem_k_index[12218] = 57105;
mem_k_index[12219] = 57108;
mem_k_index[12220] = 57110;
mem_k_index[12221] = 57113;
mem_k_index[12222] = 57115;
mem_k_index[12223] = 57118;
mem_k_index[12224] = 57120;
mem_k_index[12225] = 57123;
mem_k_index[12226] = 57125;
mem_k_index[12227] = 57128;
mem_k_index[12228] = 57130;
mem_k_index[12229] = 57133;
mem_k_index[12230] = 57135;
mem_k_index[12231] = 57138;
mem_k_index[12232] = 57140;
mem_k_index[12233] = 57143;
mem_k_index[12234] = 57145;
mem_k_index[12235] = 57148;
mem_k_index[12236] = 57150;
mem_k_index[12237] = 57153;
mem_k_index[12238] = 57155;
mem_k_index[12239] = 57158;
mem_k_index[12240] = 57160;
mem_k_index[12241] = 57163;
mem_k_index[12242] = 57165;
mem_k_index[12243] = 57168;
mem_k_index[12244] = 57170;
mem_k_index[12245] = 57173;
mem_k_index[12246] = 57176;
mem_k_index[12247] = 57178;
mem_k_index[12248] = 57181;
mem_k_index[12249] = 57183;
mem_k_index[12250] = 57186;
mem_k_index[12251] = 57188;
mem_k_index[12252] = 57191;
mem_k_index[12253] = 57193;
mem_k_index[12254] = 57196;
mem_k_index[12255] = 57198;
mem_k_index[12256] = 57201;
mem_k_index[12257] = 57203;
mem_k_index[12258] = 57206;
mem_k_index[12259] = 57208;
mem_k_index[12260] = 57211;
mem_k_index[12261] = 57213;
mem_k_index[12262] = 57216;
mem_k_index[12263] = 57218;
mem_k_index[12264] = 57221;
mem_k_index[12265] = 57223;
mem_k_index[12266] = 57226;
mem_k_index[12267] = 57228;
mem_k_index[12268] = 57231;
mem_k_index[12269] = 57233;
mem_k_index[12270] = 57236;
mem_k_index[12271] = 57238;
mem_k_index[12272] = 57241;
mem_k_index[12273] = 57243;
mem_k_index[12274] = 57246;
mem_k_index[12275] = 57248;
mem_k_index[12276] = 57251;
mem_k_index[12277] = 57253;
mem_k_index[12278] = 57256;
mem_k_index[12279] = 57258;
mem_k_index[12280] = 57261;
mem_k_index[12281] = 57263;
mem_k_index[12282] = 57266;
mem_k_index[12283] = 57268;
mem_k_index[12284] = 57271;
mem_k_index[12285] = 57273;
mem_k_index[12286] = 57276;
mem_k_index[12287] = 57278;
mem_k_index[12288] = 57600;
mem_k_index[12289] = 57602;
mem_k_index[12290] = 57605;
mem_k_index[12291] = 57607;
mem_k_index[12292] = 57610;
mem_k_index[12293] = 57612;
mem_k_index[12294] = 57615;
mem_k_index[12295] = 57617;
mem_k_index[12296] = 57620;
mem_k_index[12297] = 57622;
mem_k_index[12298] = 57625;
mem_k_index[12299] = 57627;
mem_k_index[12300] = 57630;
mem_k_index[12301] = 57632;
mem_k_index[12302] = 57635;
mem_k_index[12303] = 57637;
mem_k_index[12304] = 57640;
mem_k_index[12305] = 57642;
mem_k_index[12306] = 57645;
mem_k_index[12307] = 57647;
mem_k_index[12308] = 57650;
mem_k_index[12309] = 57652;
mem_k_index[12310] = 57655;
mem_k_index[12311] = 57657;
mem_k_index[12312] = 57660;
mem_k_index[12313] = 57662;
mem_k_index[12314] = 57665;
mem_k_index[12315] = 57667;
mem_k_index[12316] = 57670;
mem_k_index[12317] = 57672;
mem_k_index[12318] = 57675;
mem_k_index[12319] = 57677;
mem_k_index[12320] = 57680;
mem_k_index[12321] = 57682;
mem_k_index[12322] = 57685;
mem_k_index[12323] = 57687;
mem_k_index[12324] = 57690;
mem_k_index[12325] = 57692;
mem_k_index[12326] = 57695;
mem_k_index[12327] = 57697;
mem_k_index[12328] = 57700;
mem_k_index[12329] = 57702;
mem_k_index[12330] = 57705;
mem_k_index[12331] = 57708;
mem_k_index[12332] = 57710;
mem_k_index[12333] = 57713;
mem_k_index[12334] = 57715;
mem_k_index[12335] = 57718;
mem_k_index[12336] = 57720;
mem_k_index[12337] = 57723;
mem_k_index[12338] = 57725;
mem_k_index[12339] = 57728;
mem_k_index[12340] = 57730;
mem_k_index[12341] = 57733;
mem_k_index[12342] = 57735;
mem_k_index[12343] = 57738;
mem_k_index[12344] = 57740;
mem_k_index[12345] = 57743;
mem_k_index[12346] = 57745;
mem_k_index[12347] = 57748;
mem_k_index[12348] = 57750;
mem_k_index[12349] = 57753;
mem_k_index[12350] = 57755;
mem_k_index[12351] = 57758;
mem_k_index[12352] = 57760;
mem_k_index[12353] = 57763;
mem_k_index[12354] = 57765;
mem_k_index[12355] = 57768;
mem_k_index[12356] = 57770;
mem_k_index[12357] = 57773;
mem_k_index[12358] = 57775;
mem_k_index[12359] = 57778;
mem_k_index[12360] = 57780;
mem_k_index[12361] = 57783;
mem_k_index[12362] = 57785;
mem_k_index[12363] = 57788;
mem_k_index[12364] = 57790;
mem_k_index[12365] = 57793;
mem_k_index[12366] = 57795;
mem_k_index[12367] = 57798;
mem_k_index[12368] = 57800;
mem_k_index[12369] = 57803;
mem_k_index[12370] = 57805;
mem_k_index[12371] = 57808;
mem_k_index[12372] = 57810;
mem_k_index[12373] = 57813;
mem_k_index[12374] = 57816;
mem_k_index[12375] = 57818;
mem_k_index[12376] = 57821;
mem_k_index[12377] = 57823;
mem_k_index[12378] = 57826;
mem_k_index[12379] = 57828;
mem_k_index[12380] = 57831;
mem_k_index[12381] = 57833;
mem_k_index[12382] = 57836;
mem_k_index[12383] = 57838;
mem_k_index[12384] = 57841;
mem_k_index[12385] = 57843;
mem_k_index[12386] = 57846;
mem_k_index[12387] = 57848;
mem_k_index[12388] = 57851;
mem_k_index[12389] = 57853;
mem_k_index[12390] = 57856;
mem_k_index[12391] = 57858;
mem_k_index[12392] = 57861;
mem_k_index[12393] = 57863;
mem_k_index[12394] = 57866;
mem_k_index[12395] = 57868;
mem_k_index[12396] = 57871;
mem_k_index[12397] = 57873;
mem_k_index[12398] = 57876;
mem_k_index[12399] = 57878;
mem_k_index[12400] = 57881;
mem_k_index[12401] = 57883;
mem_k_index[12402] = 57886;
mem_k_index[12403] = 57888;
mem_k_index[12404] = 57891;
mem_k_index[12405] = 57893;
mem_k_index[12406] = 57896;
mem_k_index[12407] = 57898;
mem_k_index[12408] = 57901;
mem_k_index[12409] = 57903;
mem_k_index[12410] = 57906;
mem_k_index[12411] = 57908;
mem_k_index[12412] = 57911;
mem_k_index[12413] = 57913;
mem_k_index[12414] = 57916;
mem_k_index[12415] = 57918;
mem_k_index[12416] = 58240;
mem_k_index[12417] = 58242;
mem_k_index[12418] = 58245;
mem_k_index[12419] = 58247;
mem_k_index[12420] = 58250;
mem_k_index[12421] = 58252;
mem_k_index[12422] = 58255;
mem_k_index[12423] = 58257;
mem_k_index[12424] = 58260;
mem_k_index[12425] = 58262;
mem_k_index[12426] = 58265;
mem_k_index[12427] = 58267;
mem_k_index[12428] = 58270;
mem_k_index[12429] = 58272;
mem_k_index[12430] = 58275;
mem_k_index[12431] = 58277;
mem_k_index[12432] = 58280;
mem_k_index[12433] = 58282;
mem_k_index[12434] = 58285;
mem_k_index[12435] = 58287;
mem_k_index[12436] = 58290;
mem_k_index[12437] = 58292;
mem_k_index[12438] = 58295;
mem_k_index[12439] = 58297;
mem_k_index[12440] = 58300;
mem_k_index[12441] = 58302;
mem_k_index[12442] = 58305;
mem_k_index[12443] = 58307;
mem_k_index[12444] = 58310;
mem_k_index[12445] = 58312;
mem_k_index[12446] = 58315;
mem_k_index[12447] = 58317;
mem_k_index[12448] = 58320;
mem_k_index[12449] = 58322;
mem_k_index[12450] = 58325;
mem_k_index[12451] = 58327;
mem_k_index[12452] = 58330;
mem_k_index[12453] = 58332;
mem_k_index[12454] = 58335;
mem_k_index[12455] = 58337;
mem_k_index[12456] = 58340;
mem_k_index[12457] = 58342;
mem_k_index[12458] = 58345;
mem_k_index[12459] = 58348;
mem_k_index[12460] = 58350;
mem_k_index[12461] = 58353;
mem_k_index[12462] = 58355;
mem_k_index[12463] = 58358;
mem_k_index[12464] = 58360;
mem_k_index[12465] = 58363;
mem_k_index[12466] = 58365;
mem_k_index[12467] = 58368;
mem_k_index[12468] = 58370;
mem_k_index[12469] = 58373;
mem_k_index[12470] = 58375;
mem_k_index[12471] = 58378;
mem_k_index[12472] = 58380;
mem_k_index[12473] = 58383;
mem_k_index[12474] = 58385;
mem_k_index[12475] = 58388;
mem_k_index[12476] = 58390;
mem_k_index[12477] = 58393;
mem_k_index[12478] = 58395;
mem_k_index[12479] = 58398;
mem_k_index[12480] = 58400;
mem_k_index[12481] = 58403;
mem_k_index[12482] = 58405;
mem_k_index[12483] = 58408;
mem_k_index[12484] = 58410;
mem_k_index[12485] = 58413;
mem_k_index[12486] = 58415;
mem_k_index[12487] = 58418;
mem_k_index[12488] = 58420;
mem_k_index[12489] = 58423;
mem_k_index[12490] = 58425;
mem_k_index[12491] = 58428;
mem_k_index[12492] = 58430;
mem_k_index[12493] = 58433;
mem_k_index[12494] = 58435;
mem_k_index[12495] = 58438;
mem_k_index[12496] = 58440;
mem_k_index[12497] = 58443;
mem_k_index[12498] = 58445;
mem_k_index[12499] = 58448;
mem_k_index[12500] = 58450;
mem_k_index[12501] = 58453;
mem_k_index[12502] = 58456;
mem_k_index[12503] = 58458;
mem_k_index[12504] = 58461;
mem_k_index[12505] = 58463;
mem_k_index[12506] = 58466;
mem_k_index[12507] = 58468;
mem_k_index[12508] = 58471;
mem_k_index[12509] = 58473;
mem_k_index[12510] = 58476;
mem_k_index[12511] = 58478;
mem_k_index[12512] = 58481;
mem_k_index[12513] = 58483;
mem_k_index[12514] = 58486;
mem_k_index[12515] = 58488;
mem_k_index[12516] = 58491;
mem_k_index[12517] = 58493;
mem_k_index[12518] = 58496;
mem_k_index[12519] = 58498;
mem_k_index[12520] = 58501;
mem_k_index[12521] = 58503;
mem_k_index[12522] = 58506;
mem_k_index[12523] = 58508;
mem_k_index[12524] = 58511;
mem_k_index[12525] = 58513;
mem_k_index[12526] = 58516;
mem_k_index[12527] = 58518;
mem_k_index[12528] = 58521;
mem_k_index[12529] = 58523;
mem_k_index[12530] = 58526;
mem_k_index[12531] = 58528;
mem_k_index[12532] = 58531;
mem_k_index[12533] = 58533;
mem_k_index[12534] = 58536;
mem_k_index[12535] = 58538;
mem_k_index[12536] = 58541;
mem_k_index[12537] = 58543;
mem_k_index[12538] = 58546;
mem_k_index[12539] = 58548;
mem_k_index[12540] = 58551;
mem_k_index[12541] = 58553;
mem_k_index[12542] = 58556;
mem_k_index[12543] = 58558;
mem_k_index[12544] = 58880;
mem_k_index[12545] = 58882;
mem_k_index[12546] = 58885;
mem_k_index[12547] = 58887;
mem_k_index[12548] = 58890;
mem_k_index[12549] = 58892;
mem_k_index[12550] = 58895;
mem_k_index[12551] = 58897;
mem_k_index[12552] = 58900;
mem_k_index[12553] = 58902;
mem_k_index[12554] = 58905;
mem_k_index[12555] = 58907;
mem_k_index[12556] = 58910;
mem_k_index[12557] = 58912;
mem_k_index[12558] = 58915;
mem_k_index[12559] = 58917;
mem_k_index[12560] = 58920;
mem_k_index[12561] = 58922;
mem_k_index[12562] = 58925;
mem_k_index[12563] = 58927;
mem_k_index[12564] = 58930;
mem_k_index[12565] = 58932;
mem_k_index[12566] = 58935;
mem_k_index[12567] = 58937;
mem_k_index[12568] = 58940;
mem_k_index[12569] = 58942;
mem_k_index[12570] = 58945;
mem_k_index[12571] = 58947;
mem_k_index[12572] = 58950;
mem_k_index[12573] = 58952;
mem_k_index[12574] = 58955;
mem_k_index[12575] = 58957;
mem_k_index[12576] = 58960;
mem_k_index[12577] = 58962;
mem_k_index[12578] = 58965;
mem_k_index[12579] = 58967;
mem_k_index[12580] = 58970;
mem_k_index[12581] = 58972;
mem_k_index[12582] = 58975;
mem_k_index[12583] = 58977;
mem_k_index[12584] = 58980;
mem_k_index[12585] = 58982;
mem_k_index[12586] = 58985;
mem_k_index[12587] = 58988;
mem_k_index[12588] = 58990;
mem_k_index[12589] = 58993;
mem_k_index[12590] = 58995;
mem_k_index[12591] = 58998;
mem_k_index[12592] = 59000;
mem_k_index[12593] = 59003;
mem_k_index[12594] = 59005;
mem_k_index[12595] = 59008;
mem_k_index[12596] = 59010;
mem_k_index[12597] = 59013;
mem_k_index[12598] = 59015;
mem_k_index[12599] = 59018;
mem_k_index[12600] = 59020;
mem_k_index[12601] = 59023;
mem_k_index[12602] = 59025;
mem_k_index[12603] = 59028;
mem_k_index[12604] = 59030;
mem_k_index[12605] = 59033;
mem_k_index[12606] = 59035;
mem_k_index[12607] = 59038;
mem_k_index[12608] = 59040;
mem_k_index[12609] = 59043;
mem_k_index[12610] = 59045;
mem_k_index[12611] = 59048;
mem_k_index[12612] = 59050;
mem_k_index[12613] = 59053;
mem_k_index[12614] = 59055;
mem_k_index[12615] = 59058;
mem_k_index[12616] = 59060;
mem_k_index[12617] = 59063;
mem_k_index[12618] = 59065;
mem_k_index[12619] = 59068;
mem_k_index[12620] = 59070;
mem_k_index[12621] = 59073;
mem_k_index[12622] = 59075;
mem_k_index[12623] = 59078;
mem_k_index[12624] = 59080;
mem_k_index[12625] = 59083;
mem_k_index[12626] = 59085;
mem_k_index[12627] = 59088;
mem_k_index[12628] = 59090;
mem_k_index[12629] = 59093;
mem_k_index[12630] = 59096;
mem_k_index[12631] = 59098;
mem_k_index[12632] = 59101;
mem_k_index[12633] = 59103;
mem_k_index[12634] = 59106;
mem_k_index[12635] = 59108;
mem_k_index[12636] = 59111;
mem_k_index[12637] = 59113;
mem_k_index[12638] = 59116;
mem_k_index[12639] = 59118;
mem_k_index[12640] = 59121;
mem_k_index[12641] = 59123;
mem_k_index[12642] = 59126;
mem_k_index[12643] = 59128;
mem_k_index[12644] = 59131;
mem_k_index[12645] = 59133;
mem_k_index[12646] = 59136;
mem_k_index[12647] = 59138;
mem_k_index[12648] = 59141;
mem_k_index[12649] = 59143;
mem_k_index[12650] = 59146;
mem_k_index[12651] = 59148;
mem_k_index[12652] = 59151;
mem_k_index[12653] = 59153;
mem_k_index[12654] = 59156;
mem_k_index[12655] = 59158;
mem_k_index[12656] = 59161;
mem_k_index[12657] = 59163;
mem_k_index[12658] = 59166;
mem_k_index[12659] = 59168;
mem_k_index[12660] = 59171;
mem_k_index[12661] = 59173;
mem_k_index[12662] = 59176;
mem_k_index[12663] = 59178;
mem_k_index[12664] = 59181;
mem_k_index[12665] = 59183;
mem_k_index[12666] = 59186;
mem_k_index[12667] = 59188;
mem_k_index[12668] = 59191;
mem_k_index[12669] = 59193;
mem_k_index[12670] = 59196;
mem_k_index[12671] = 59198;
mem_k_index[12672] = 59520;
mem_k_index[12673] = 59522;
mem_k_index[12674] = 59525;
mem_k_index[12675] = 59527;
mem_k_index[12676] = 59530;
mem_k_index[12677] = 59532;
mem_k_index[12678] = 59535;
mem_k_index[12679] = 59537;
mem_k_index[12680] = 59540;
mem_k_index[12681] = 59542;
mem_k_index[12682] = 59545;
mem_k_index[12683] = 59547;
mem_k_index[12684] = 59550;
mem_k_index[12685] = 59552;
mem_k_index[12686] = 59555;
mem_k_index[12687] = 59557;
mem_k_index[12688] = 59560;
mem_k_index[12689] = 59562;
mem_k_index[12690] = 59565;
mem_k_index[12691] = 59567;
mem_k_index[12692] = 59570;
mem_k_index[12693] = 59572;
mem_k_index[12694] = 59575;
mem_k_index[12695] = 59577;
mem_k_index[12696] = 59580;
mem_k_index[12697] = 59582;
mem_k_index[12698] = 59585;
mem_k_index[12699] = 59587;
mem_k_index[12700] = 59590;
mem_k_index[12701] = 59592;
mem_k_index[12702] = 59595;
mem_k_index[12703] = 59597;
mem_k_index[12704] = 59600;
mem_k_index[12705] = 59602;
mem_k_index[12706] = 59605;
mem_k_index[12707] = 59607;
mem_k_index[12708] = 59610;
mem_k_index[12709] = 59612;
mem_k_index[12710] = 59615;
mem_k_index[12711] = 59617;
mem_k_index[12712] = 59620;
mem_k_index[12713] = 59622;
mem_k_index[12714] = 59625;
mem_k_index[12715] = 59628;
mem_k_index[12716] = 59630;
mem_k_index[12717] = 59633;
mem_k_index[12718] = 59635;
mem_k_index[12719] = 59638;
mem_k_index[12720] = 59640;
mem_k_index[12721] = 59643;
mem_k_index[12722] = 59645;
mem_k_index[12723] = 59648;
mem_k_index[12724] = 59650;
mem_k_index[12725] = 59653;
mem_k_index[12726] = 59655;
mem_k_index[12727] = 59658;
mem_k_index[12728] = 59660;
mem_k_index[12729] = 59663;
mem_k_index[12730] = 59665;
mem_k_index[12731] = 59668;
mem_k_index[12732] = 59670;
mem_k_index[12733] = 59673;
mem_k_index[12734] = 59675;
mem_k_index[12735] = 59678;
mem_k_index[12736] = 59680;
mem_k_index[12737] = 59683;
mem_k_index[12738] = 59685;
mem_k_index[12739] = 59688;
mem_k_index[12740] = 59690;
mem_k_index[12741] = 59693;
mem_k_index[12742] = 59695;
mem_k_index[12743] = 59698;
mem_k_index[12744] = 59700;
mem_k_index[12745] = 59703;
mem_k_index[12746] = 59705;
mem_k_index[12747] = 59708;
mem_k_index[12748] = 59710;
mem_k_index[12749] = 59713;
mem_k_index[12750] = 59715;
mem_k_index[12751] = 59718;
mem_k_index[12752] = 59720;
mem_k_index[12753] = 59723;
mem_k_index[12754] = 59725;
mem_k_index[12755] = 59728;
mem_k_index[12756] = 59730;
mem_k_index[12757] = 59733;
mem_k_index[12758] = 59736;
mem_k_index[12759] = 59738;
mem_k_index[12760] = 59741;
mem_k_index[12761] = 59743;
mem_k_index[12762] = 59746;
mem_k_index[12763] = 59748;
mem_k_index[12764] = 59751;
mem_k_index[12765] = 59753;
mem_k_index[12766] = 59756;
mem_k_index[12767] = 59758;
mem_k_index[12768] = 59761;
mem_k_index[12769] = 59763;
mem_k_index[12770] = 59766;
mem_k_index[12771] = 59768;
mem_k_index[12772] = 59771;
mem_k_index[12773] = 59773;
mem_k_index[12774] = 59776;
mem_k_index[12775] = 59778;
mem_k_index[12776] = 59781;
mem_k_index[12777] = 59783;
mem_k_index[12778] = 59786;
mem_k_index[12779] = 59788;
mem_k_index[12780] = 59791;
mem_k_index[12781] = 59793;
mem_k_index[12782] = 59796;
mem_k_index[12783] = 59798;
mem_k_index[12784] = 59801;
mem_k_index[12785] = 59803;
mem_k_index[12786] = 59806;
mem_k_index[12787] = 59808;
mem_k_index[12788] = 59811;
mem_k_index[12789] = 59813;
mem_k_index[12790] = 59816;
mem_k_index[12791] = 59818;
mem_k_index[12792] = 59821;
mem_k_index[12793] = 59823;
mem_k_index[12794] = 59826;
mem_k_index[12795] = 59828;
mem_k_index[12796] = 59831;
mem_k_index[12797] = 59833;
mem_k_index[12798] = 59836;
mem_k_index[12799] = 59838;
mem_k_index[12800] = 60160;
mem_k_index[12801] = 60162;
mem_k_index[12802] = 60165;
mem_k_index[12803] = 60167;
mem_k_index[12804] = 60170;
mem_k_index[12805] = 60172;
mem_k_index[12806] = 60175;
mem_k_index[12807] = 60177;
mem_k_index[12808] = 60180;
mem_k_index[12809] = 60182;
mem_k_index[12810] = 60185;
mem_k_index[12811] = 60187;
mem_k_index[12812] = 60190;
mem_k_index[12813] = 60192;
mem_k_index[12814] = 60195;
mem_k_index[12815] = 60197;
mem_k_index[12816] = 60200;
mem_k_index[12817] = 60202;
mem_k_index[12818] = 60205;
mem_k_index[12819] = 60207;
mem_k_index[12820] = 60210;
mem_k_index[12821] = 60212;
mem_k_index[12822] = 60215;
mem_k_index[12823] = 60217;
mem_k_index[12824] = 60220;
mem_k_index[12825] = 60222;
mem_k_index[12826] = 60225;
mem_k_index[12827] = 60227;
mem_k_index[12828] = 60230;
mem_k_index[12829] = 60232;
mem_k_index[12830] = 60235;
mem_k_index[12831] = 60237;
mem_k_index[12832] = 60240;
mem_k_index[12833] = 60242;
mem_k_index[12834] = 60245;
mem_k_index[12835] = 60247;
mem_k_index[12836] = 60250;
mem_k_index[12837] = 60252;
mem_k_index[12838] = 60255;
mem_k_index[12839] = 60257;
mem_k_index[12840] = 60260;
mem_k_index[12841] = 60262;
mem_k_index[12842] = 60265;
mem_k_index[12843] = 60268;
mem_k_index[12844] = 60270;
mem_k_index[12845] = 60273;
mem_k_index[12846] = 60275;
mem_k_index[12847] = 60278;
mem_k_index[12848] = 60280;
mem_k_index[12849] = 60283;
mem_k_index[12850] = 60285;
mem_k_index[12851] = 60288;
mem_k_index[12852] = 60290;
mem_k_index[12853] = 60293;
mem_k_index[12854] = 60295;
mem_k_index[12855] = 60298;
mem_k_index[12856] = 60300;
mem_k_index[12857] = 60303;
mem_k_index[12858] = 60305;
mem_k_index[12859] = 60308;
mem_k_index[12860] = 60310;
mem_k_index[12861] = 60313;
mem_k_index[12862] = 60315;
mem_k_index[12863] = 60318;
mem_k_index[12864] = 60320;
mem_k_index[12865] = 60323;
mem_k_index[12866] = 60325;
mem_k_index[12867] = 60328;
mem_k_index[12868] = 60330;
mem_k_index[12869] = 60333;
mem_k_index[12870] = 60335;
mem_k_index[12871] = 60338;
mem_k_index[12872] = 60340;
mem_k_index[12873] = 60343;
mem_k_index[12874] = 60345;
mem_k_index[12875] = 60348;
mem_k_index[12876] = 60350;
mem_k_index[12877] = 60353;
mem_k_index[12878] = 60355;
mem_k_index[12879] = 60358;
mem_k_index[12880] = 60360;
mem_k_index[12881] = 60363;
mem_k_index[12882] = 60365;
mem_k_index[12883] = 60368;
mem_k_index[12884] = 60370;
mem_k_index[12885] = 60373;
mem_k_index[12886] = 60376;
mem_k_index[12887] = 60378;
mem_k_index[12888] = 60381;
mem_k_index[12889] = 60383;
mem_k_index[12890] = 60386;
mem_k_index[12891] = 60388;
mem_k_index[12892] = 60391;
mem_k_index[12893] = 60393;
mem_k_index[12894] = 60396;
mem_k_index[12895] = 60398;
mem_k_index[12896] = 60401;
mem_k_index[12897] = 60403;
mem_k_index[12898] = 60406;
mem_k_index[12899] = 60408;
mem_k_index[12900] = 60411;
mem_k_index[12901] = 60413;
mem_k_index[12902] = 60416;
mem_k_index[12903] = 60418;
mem_k_index[12904] = 60421;
mem_k_index[12905] = 60423;
mem_k_index[12906] = 60426;
mem_k_index[12907] = 60428;
mem_k_index[12908] = 60431;
mem_k_index[12909] = 60433;
mem_k_index[12910] = 60436;
mem_k_index[12911] = 60438;
mem_k_index[12912] = 60441;
mem_k_index[12913] = 60443;
mem_k_index[12914] = 60446;
mem_k_index[12915] = 60448;
mem_k_index[12916] = 60451;
mem_k_index[12917] = 60453;
mem_k_index[12918] = 60456;
mem_k_index[12919] = 60458;
mem_k_index[12920] = 60461;
mem_k_index[12921] = 60463;
mem_k_index[12922] = 60466;
mem_k_index[12923] = 60468;
mem_k_index[12924] = 60471;
mem_k_index[12925] = 60473;
mem_k_index[12926] = 60476;
mem_k_index[12927] = 60478;
mem_k_index[12928] = 60800;
mem_k_index[12929] = 60802;
mem_k_index[12930] = 60805;
mem_k_index[12931] = 60807;
mem_k_index[12932] = 60810;
mem_k_index[12933] = 60812;
mem_k_index[12934] = 60815;
mem_k_index[12935] = 60817;
mem_k_index[12936] = 60820;
mem_k_index[12937] = 60822;
mem_k_index[12938] = 60825;
mem_k_index[12939] = 60827;
mem_k_index[12940] = 60830;
mem_k_index[12941] = 60832;
mem_k_index[12942] = 60835;
mem_k_index[12943] = 60837;
mem_k_index[12944] = 60840;
mem_k_index[12945] = 60842;
mem_k_index[12946] = 60845;
mem_k_index[12947] = 60847;
mem_k_index[12948] = 60850;
mem_k_index[12949] = 60852;
mem_k_index[12950] = 60855;
mem_k_index[12951] = 60857;
mem_k_index[12952] = 60860;
mem_k_index[12953] = 60862;
mem_k_index[12954] = 60865;
mem_k_index[12955] = 60867;
mem_k_index[12956] = 60870;
mem_k_index[12957] = 60872;
mem_k_index[12958] = 60875;
mem_k_index[12959] = 60877;
mem_k_index[12960] = 60880;
mem_k_index[12961] = 60882;
mem_k_index[12962] = 60885;
mem_k_index[12963] = 60887;
mem_k_index[12964] = 60890;
mem_k_index[12965] = 60892;
mem_k_index[12966] = 60895;
mem_k_index[12967] = 60897;
mem_k_index[12968] = 60900;
mem_k_index[12969] = 60902;
mem_k_index[12970] = 60905;
mem_k_index[12971] = 60908;
mem_k_index[12972] = 60910;
mem_k_index[12973] = 60913;
mem_k_index[12974] = 60915;
mem_k_index[12975] = 60918;
mem_k_index[12976] = 60920;
mem_k_index[12977] = 60923;
mem_k_index[12978] = 60925;
mem_k_index[12979] = 60928;
mem_k_index[12980] = 60930;
mem_k_index[12981] = 60933;
mem_k_index[12982] = 60935;
mem_k_index[12983] = 60938;
mem_k_index[12984] = 60940;
mem_k_index[12985] = 60943;
mem_k_index[12986] = 60945;
mem_k_index[12987] = 60948;
mem_k_index[12988] = 60950;
mem_k_index[12989] = 60953;
mem_k_index[12990] = 60955;
mem_k_index[12991] = 60958;
mem_k_index[12992] = 60960;
mem_k_index[12993] = 60963;
mem_k_index[12994] = 60965;
mem_k_index[12995] = 60968;
mem_k_index[12996] = 60970;
mem_k_index[12997] = 60973;
mem_k_index[12998] = 60975;
mem_k_index[12999] = 60978;
mem_k_index[13000] = 60980;
mem_k_index[13001] = 60983;
mem_k_index[13002] = 60985;
mem_k_index[13003] = 60988;
mem_k_index[13004] = 60990;
mem_k_index[13005] = 60993;
mem_k_index[13006] = 60995;
mem_k_index[13007] = 60998;
mem_k_index[13008] = 61000;
mem_k_index[13009] = 61003;
mem_k_index[13010] = 61005;
mem_k_index[13011] = 61008;
mem_k_index[13012] = 61010;
mem_k_index[13013] = 61013;
mem_k_index[13014] = 61016;
mem_k_index[13015] = 61018;
mem_k_index[13016] = 61021;
mem_k_index[13017] = 61023;
mem_k_index[13018] = 61026;
mem_k_index[13019] = 61028;
mem_k_index[13020] = 61031;
mem_k_index[13021] = 61033;
mem_k_index[13022] = 61036;
mem_k_index[13023] = 61038;
mem_k_index[13024] = 61041;
mem_k_index[13025] = 61043;
mem_k_index[13026] = 61046;
mem_k_index[13027] = 61048;
mem_k_index[13028] = 61051;
mem_k_index[13029] = 61053;
mem_k_index[13030] = 61056;
mem_k_index[13031] = 61058;
mem_k_index[13032] = 61061;
mem_k_index[13033] = 61063;
mem_k_index[13034] = 61066;
mem_k_index[13035] = 61068;
mem_k_index[13036] = 61071;
mem_k_index[13037] = 61073;
mem_k_index[13038] = 61076;
mem_k_index[13039] = 61078;
mem_k_index[13040] = 61081;
mem_k_index[13041] = 61083;
mem_k_index[13042] = 61086;
mem_k_index[13043] = 61088;
mem_k_index[13044] = 61091;
mem_k_index[13045] = 61093;
mem_k_index[13046] = 61096;
mem_k_index[13047] = 61098;
mem_k_index[13048] = 61101;
mem_k_index[13049] = 61103;
mem_k_index[13050] = 61106;
mem_k_index[13051] = 61108;
mem_k_index[13052] = 61111;
mem_k_index[13053] = 61113;
mem_k_index[13054] = 61116;
mem_k_index[13055] = 61118;
mem_k_index[13056] = 61120;
mem_k_index[13057] = 61122;
mem_k_index[13058] = 61125;
mem_k_index[13059] = 61127;
mem_k_index[13060] = 61130;
mem_k_index[13061] = 61132;
mem_k_index[13062] = 61135;
mem_k_index[13063] = 61137;
mem_k_index[13064] = 61140;
mem_k_index[13065] = 61142;
mem_k_index[13066] = 61145;
mem_k_index[13067] = 61147;
mem_k_index[13068] = 61150;
mem_k_index[13069] = 61152;
mem_k_index[13070] = 61155;
mem_k_index[13071] = 61157;
mem_k_index[13072] = 61160;
mem_k_index[13073] = 61162;
mem_k_index[13074] = 61165;
mem_k_index[13075] = 61167;
mem_k_index[13076] = 61170;
mem_k_index[13077] = 61172;
mem_k_index[13078] = 61175;
mem_k_index[13079] = 61177;
mem_k_index[13080] = 61180;
mem_k_index[13081] = 61182;
mem_k_index[13082] = 61185;
mem_k_index[13083] = 61187;
mem_k_index[13084] = 61190;
mem_k_index[13085] = 61192;
mem_k_index[13086] = 61195;
mem_k_index[13087] = 61197;
mem_k_index[13088] = 61200;
mem_k_index[13089] = 61202;
mem_k_index[13090] = 61205;
mem_k_index[13091] = 61207;
mem_k_index[13092] = 61210;
mem_k_index[13093] = 61212;
mem_k_index[13094] = 61215;
mem_k_index[13095] = 61217;
mem_k_index[13096] = 61220;
mem_k_index[13097] = 61222;
mem_k_index[13098] = 61225;
mem_k_index[13099] = 61228;
mem_k_index[13100] = 61230;
mem_k_index[13101] = 61233;
mem_k_index[13102] = 61235;
mem_k_index[13103] = 61238;
mem_k_index[13104] = 61240;
mem_k_index[13105] = 61243;
mem_k_index[13106] = 61245;
mem_k_index[13107] = 61248;
mem_k_index[13108] = 61250;
mem_k_index[13109] = 61253;
mem_k_index[13110] = 61255;
mem_k_index[13111] = 61258;
mem_k_index[13112] = 61260;
mem_k_index[13113] = 61263;
mem_k_index[13114] = 61265;
mem_k_index[13115] = 61268;
mem_k_index[13116] = 61270;
mem_k_index[13117] = 61273;
mem_k_index[13118] = 61275;
mem_k_index[13119] = 61278;
mem_k_index[13120] = 61280;
mem_k_index[13121] = 61283;
mem_k_index[13122] = 61285;
mem_k_index[13123] = 61288;
mem_k_index[13124] = 61290;
mem_k_index[13125] = 61293;
mem_k_index[13126] = 61295;
mem_k_index[13127] = 61298;
mem_k_index[13128] = 61300;
mem_k_index[13129] = 61303;
mem_k_index[13130] = 61305;
mem_k_index[13131] = 61308;
mem_k_index[13132] = 61310;
mem_k_index[13133] = 61313;
mem_k_index[13134] = 61315;
mem_k_index[13135] = 61318;
mem_k_index[13136] = 61320;
mem_k_index[13137] = 61323;
mem_k_index[13138] = 61325;
mem_k_index[13139] = 61328;
mem_k_index[13140] = 61330;
mem_k_index[13141] = 61333;
mem_k_index[13142] = 61336;
mem_k_index[13143] = 61338;
mem_k_index[13144] = 61341;
mem_k_index[13145] = 61343;
mem_k_index[13146] = 61346;
mem_k_index[13147] = 61348;
mem_k_index[13148] = 61351;
mem_k_index[13149] = 61353;
mem_k_index[13150] = 61356;
mem_k_index[13151] = 61358;
mem_k_index[13152] = 61361;
mem_k_index[13153] = 61363;
mem_k_index[13154] = 61366;
mem_k_index[13155] = 61368;
mem_k_index[13156] = 61371;
mem_k_index[13157] = 61373;
mem_k_index[13158] = 61376;
mem_k_index[13159] = 61378;
mem_k_index[13160] = 61381;
mem_k_index[13161] = 61383;
mem_k_index[13162] = 61386;
mem_k_index[13163] = 61388;
mem_k_index[13164] = 61391;
mem_k_index[13165] = 61393;
mem_k_index[13166] = 61396;
mem_k_index[13167] = 61398;
mem_k_index[13168] = 61401;
mem_k_index[13169] = 61403;
mem_k_index[13170] = 61406;
mem_k_index[13171] = 61408;
mem_k_index[13172] = 61411;
mem_k_index[13173] = 61413;
mem_k_index[13174] = 61416;
mem_k_index[13175] = 61418;
mem_k_index[13176] = 61421;
mem_k_index[13177] = 61423;
mem_k_index[13178] = 61426;
mem_k_index[13179] = 61428;
mem_k_index[13180] = 61431;
mem_k_index[13181] = 61433;
mem_k_index[13182] = 61436;
mem_k_index[13183] = 61438;
mem_k_index[13184] = 61760;
mem_k_index[13185] = 61762;
mem_k_index[13186] = 61765;
mem_k_index[13187] = 61767;
mem_k_index[13188] = 61770;
mem_k_index[13189] = 61772;
mem_k_index[13190] = 61775;
mem_k_index[13191] = 61777;
mem_k_index[13192] = 61780;
mem_k_index[13193] = 61782;
mem_k_index[13194] = 61785;
mem_k_index[13195] = 61787;
mem_k_index[13196] = 61790;
mem_k_index[13197] = 61792;
mem_k_index[13198] = 61795;
mem_k_index[13199] = 61797;
mem_k_index[13200] = 61800;
mem_k_index[13201] = 61802;
mem_k_index[13202] = 61805;
mem_k_index[13203] = 61807;
mem_k_index[13204] = 61810;
mem_k_index[13205] = 61812;
mem_k_index[13206] = 61815;
mem_k_index[13207] = 61817;
mem_k_index[13208] = 61820;
mem_k_index[13209] = 61822;
mem_k_index[13210] = 61825;
mem_k_index[13211] = 61827;
mem_k_index[13212] = 61830;
mem_k_index[13213] = 61832;
mem_k_index[13214] = 61835;
mem_k_index[13215] = 61837;
mem_k_index[13216] = 61840;
mem_k_index[13217] = 61842;
mem_k_index[13218] = 61845;
mem_k_index[13219] = 61847;
mem_k_index[13220] = 61850;
mem_k_index[13221] = 61852;
mem_k_index[13222] = 61855;
mem_k_index[13223] = 61857;
mem_k_index[13224] = 61860;
mem_k_index[13225] = 61862;
mem_k_index[13226] = 61865;
mem_k_index[13227] = 61868;
mem_k_index[13228] = 61870;
mem_k_index[13229] = 61873;
mem_k_index[13230] = 61875;
mem_k_index[13231] = 61878;
mem_k_index[13232] = 61880;
mem_k_index[13233] = 61883;
mem_k_index[13234] = 61885;
mem_k_index[13235] = 61888;
mem_k_index[13236] = 61890;
mem_k_index[13237] = 61893;
mem_k_index[13238] = 61895;
mem_k_index[13239] = 61898;
mem_k_index[13240] = 61900;
mem_k_index[13241] = 61903;
mem_k_index[13242] = 61905;
mem_k_index[13243] = 61908;
mem_k_index[13244] = 61910;
mem_k_index[13245] = 61913;
mem_k_index[13246] = 61915;
mem_k_index[13247] = 61918;
mem_k_index[13248] = 61920;
mem_k_index[13249] = 61923;
mem_k_index[13250] = 61925;
mem_k_index[13251] = 61928;
mem_k_index[13252] = 61930;
mem_k_index[13253] = 61933;
mem_k_index[13254] = 61935;
mem_k_index[13255] = 61938;
mem_k_index[13256] = 61940;
mem_k_index[13257] = 61943;
mem_k_index[13258] = 61945;
mem_k_index[13259] = 61948;
mem_k_index[13260] = 61950;
mem_k_index[13261] = 61953;
mem_k_index[13262] = 61955;
mem_k_index[13263] = 61958;
mem_k_index[13264] = 61960;
mem_k_index[13265] = 61963;
mem_k_index[13266] = 61965;
mem_k_index[13267] = 61968;
mem_k_index[13268] = 61970;
mem_k_index[13269] = 61973;
mem_k_index[13270] = 61976;
mem_k_index[13271] = 61978;
mem_k_index[13272] = 61981;
mem_k_index[13273] = 61983;
mem_k_index[13274] = 61986;
mem_k_index[13275] = 61988;
mem_k_index[13276] = 61991;
mem_k_index[13277] = 61993;
mem_k_index[13278] = 61996;
mem_k_index[13279] = 61998;
mem_k_index[13280] = 62001;
mem_k_index[13281] = 62003;
mem_k_index[13282] = 62006;
mem_k_index[13283] = 62008;
mem_k_index[13284] = 62011;
mem_k_index[13285] = 62013;
mem_k_index[13286] = 62016;
mem_k_index[13287] = 62018;
mem_k_index[13288] = 62021;
mem_k_index[13289] = 62023;
mem_k_index[13290] = 62026;
mem_k_index[13291] = 62028;
mem_k_index[13292] = 62031;
mem_k_index[13293] = 62033;
mem_k_index[13294] = 62036;
mem_k_index[13295] = 62038;
mem_k_index[13296] = 62041;
mem_k_index[13297] = 62043;
mem_k_index[13298] = 62046;
mem_k_index[13299] = 62048;
mem_k_index[13300] = 62051;
mem_k_index[13301] = 62053;
mem_k_index[13302] = 62056;
mem_k_index[13303] = 62058;
mem_k_index[13304] = 62061;
mem_k_index[13305] = 62063;
mem_k_index[13306] = 62066;
mem_k_index[13307] = 62068;
mem_k_index[13308] = 62071;
mem_k_index[13309] = 62073;
mem_k_index[13310] = 62076;
mem_k_index[13311] = 62078;
mem_k_index[13312] = 62400;
mem_k_index[13313] = 62402;
mem_k_index[13314] = 62405;
mem_k_index[13315] = 62407;
mem_k_index[13316] = 62410;
mem_k_index[13317] = 62412;
mem_k_index[13318] = 62415;
mem_k_index[13319] = 62417;
mem_k_index[13320] = 62420;
mem_k_index[13321] = 62422;
mem_k_index[13322] = 62425;
mem_k_index[13323] = 62427;
mem_k_index[13324] = 62430;
mem_k_index[13325] = 62432;
mem_k_index[13326] = 62435;
mem_k_index[13327] = 62437;
mem_k_index[13328] = 62440;
mem_k_index[13329] = 62442;
mem_k_index[13330] = 62445;
mem_k_index[13331] = 62447;
mem_k_index[13332] = 62450;
mem_k_index[13333] = 62452;
mem_k_index[13334] = 62455;
mem_k_index[13335] = 62457;
mem_k_index[13336] = 62460;
mem_k_index[13337] = 62462;
mem_k_index[13338] = 62465;
mem_k_index[13339] = 62467;
mem_k_index[13340] = 62470;
mem_k_index[13341] = 62472;
mem_k_index[13342] = 62475;
mem_k_index[13343] = 62477;
mem_k_index[13344] = 62480;
mem_k_index[13345] = 62482;
mem_k_index[13346] = 62485;
mem_k_index[13347] = 62487;
mem_k_index[13348] = 62490;
mem_k_index[13349] = 62492;
mem_k_index[13350] = 62495;
mem_k_index[13351] = 62497;
mem_k_index[13352] = 62500;
mem_k_index[13353] = 62502;
mem_k_index[13354] = 62505;
mem_k_index[13355] = 62508;
mem_k_index[13356] = 62510;
mem_k_index[13357] = 62513;
mem_k_index[13358] = 62515;
mem_k_index[13359] = 62518;
mem_k_index[13360] = 62520;
mem_k_index[13361] = 62523;
mem_k_index[13362] = 62525;
mem_k_index[13363] = 62528;
mem_k_index[13364] = 62530;
mem_k_index[13365] = 62533;
mem_k_index[13366] = 62535;
mem_k_index[13367] = 62538;
mem_k_index[13368] = 62540;
mem_k_index[13369] = 62543;
mem_k_index[13370] = 62545;
mem_k_index[13371] = 62548;
mem_k_index[13372] = 62550;
mem_k_index[13373] = 62553;
mem_k_index[13374] = 62555;
mem_k_index[13375] = 62558;
mem_k_index[13376] = 62560;
mem_k_index[13377] = 62563;
mem_k_index[13378] = 62565;
mem_k_index[13379] = 62568;
mem_k_index[13380] = 62570;
mem_k_index[13381] = 62573;
mem_k_index[13382] = 62575;
mem_k_index[13383] = 62578;
mem_k_index[13384] = 62580;
mem_k_index[13385] = 62583;
mem_k_index[13386] = 62585;
mem_k_index[13387] = 62588;
mem_k_index[13388] = 62590;
mem_k_index[13389] = 62593;
mem_k_index[13390] = 62595;
mem_k_index[13391] = 62598;
mem_k_index[13392] = 62600;
mem_k_index[13393] = 62603;
mem_k_index[13394] = 62605;
mem_k_index[13395] = 62608;
mem_k_index[13396] = 62610;
mem_k_index[13397] = 62613;
mem_k_index[13398] = 62616;
mem_k_index[13399] = 62618;
mem_k_index[13400] = 62621;
mem_k_index[13401] = 62623;
mem_k_index[13402] = 62626;
mem_k_index[13403] = 62628;
mem_k_index[13404] = 62631;
mem_k_index[13405] = 62633;
mem_k_index[13406] = 62636;
mem_k_index[13407] = 62638;
mem_k_index[13408] = 62641;
mem_k_index[13409] = 62643;
mem_k_index[13410] = 62646;
mem_k_index[13411] = 62648;
mem_k_index[13412] = 62651;
mem_k_index[13413] = 62653;
mem_k_index[13414] = 62656;
mem_k_index[13415] = 62658;
mem_k_index[13416] = 62661;
mem_k_index[13417] = 62663;
mem_k_index[13418] = 62666;
mem_k_index[13419] = 62668;
mem_k_index[13420] = 62671;
mem_k_index[13421] = 62673;
mem_k_index[13422] = 62676;
mem_k_index[13423] = 62678;
mem_k_index[13424] = 62681;
mem_k_index[13425] = 62683;
mem_k_index[13426] = 62686;
mem_k_index[13427] = 62688;
mem_k_index[13428] = 62691;
mem_k_index[13429] = 62693;
mem_k_index[13430] = 62696;
mem_k_index[13431] = 62698;
mem_k_index[13432] = 62701;
mem_k_index[13433] = 62703;
mem_k_index[13434] = 62706;
mem_k_index[13435] = 62708;
mem_k_index[13436] = 62711;
mem_k_index[13437] = 62713;
mem_k_index[13438] = 62716;
mem_k_index[13439] = 62718;
mem_k_index[13440] = 63040;
mem_k_index[13441] = 63042;
mem_k_index[13442] = 63045;
mem_k_index[13443] = 63047;
mem_k_index[13444] = 63050;
mem_k_index[13445] = 63052;
mem_k_index[13446] = 63055;
mem_k_index[13447] = 63057;
mem_k_index[13448] = 63060;
mem_k_index[13449] = 63062;
mem_k_index[13450] = 63065;
mem_k_index[13451] = 63067;
mem_k_index[13452] = 63070;
mem_k_index[13453] = 63072;
mem_k_index[13454] = 63075;
mem_k_index[13455] = 63077;
mem_k_index[13456] = 63080;
mem_k_index[13457] = 63082;
mem_k_index[13458] = 63085;
mem_k_index[13459] = 63087;
mem_k_index[13460] = 63090;
mem_k_index[13461] = 63092;
mem_k_index[13462] = 63095;
mem_k_index[13463] = 63097;
mem_k_index[13464] = 63100;
mem_k_index[13465] = 63102;
mem_k_index[13466] = 63105;
mem_k_index[13467] = 63107;
mem_k_index[13468] = 63110;
mem_k_index[13469] = 63112;
mem_k_index[13470] = 63115;
mem_k_index[13471] = 63117;
mem_k_index[13472] = 63120;
mem_k_index[13473] = 63122;
mem_k_index[13474] = 63125;
mem_k_index[13475] = 63127;
mem_k_index[13476] = 63130;
mem_k_index[13477] = 63132;
mem_k_index[13478] = 63135;
mem_k_index[13479] = 63137;
mem_k_index[13480] = 63140;
mem_k_index[13481] = 63142;
mem_k_index[13482] = 63145;
mem_k_index[13483] = 63148;
mem_k_index[13484] = 63150;
mem_k_index[13485] = 63153;
mem_k_index[13486] = 63155;
mem_k_index[13487] = 63158;
mem_k_index[13488] = 63160;
mem_k_index[13489] = 63163;
mem_k_index[13490] = 63165;
mem_k_index[13491] = 63168;
mem_k_index[13492] = 63170;
mem_k_index[13493] = 63173;
mem_k_index[13494] = 63175;
mem_k_index[13495] = 63178;
mem_k_index[13496] = 63180;
mem_k_index[13497] = 63183;
mem_k_index[13498] = 63185;
mem_k_index[13499] = 63188;
mem_k_index[13500] = 63190;
mem_k_index[13501] = 63193;
mem_k_index[13502] = 63195;
mem_k_index[13503] = 63198;
mem_k_index[13504] = 63200;
mem_k_index[13505] = 63203;
mem_k_index[13506] = 63205;
mem_k_index[13507] = 63208;
mem_k_index[13508] = 63210;
mem_k_index[13509] = 63213;
mem_k_index[13510] = 63215;
mem_k_index[13511] = 63218;
mem_k_index[13512] = 63220;
mem_k_index[13513] = 63223;
mem_k_index[13514] = 63225;
mem_k_index[13515] = 63228;
mem_k_index[13516] = 63230;
mem_k_index[13517] = 63233;
mem_k_index[13518] = 63235;
mem_k_index[13519] = 63238;
mem_k_index[13520] = 63240;
mem_k_index[13521] = 63243;
mem_k_index[13522] = 63245;
mem_k_index[13523] = 63248;
mem_k_index[13524] = 63250;
mem_k_index[13525] = 63253;
mem_k_index[13526] = 63256;
mem_k_index[13527] = 63258;
mem_k_index[13528] = 63261;
mem_k_index[13529] = 63263;
mem_k_index[13530] = 63266;
mem_k_index[13531] = 63268;
mem_k_index[13532] = 63271;
mem_k_index[13533] = 63273;
mem_k_index[13534] = 63276;
mem_k_index[13535] = 63278;
mem_k_index[13536] = 63281;
mem_k_index[13537] = 63283;
mem_k_index[13538] = 63286;
mem_k_index[13539] = 63288;
mem_k_index[13540] = 63291;
mem_k_index[13541] = 63293;
mem_k_index[13542] = 63296;
mem_k_index[13543] = 63298;
mem_k_index[13544] = 63301;
mem_k_index[13545] = 63303;
mem_k_index[13546] = 63306;
mem_k_index[13547] = 63308;
mem_k_index[13548] = 63311;
mem_k_index[13549] = 63313;
mem_k_index[13550] = 63316;
mem_k_index[13551] = 63318;
mem_k_index[13552] = 63321;
mem_k_index[13553] = 63323;
mem_k_index[13554] = 63326;
mem_k_index[13555] = 63328;
mem_k_index[13556] = 63331;
mem_k_index[13557] = 63333;
mem_k_index[13558] = 63336;
mem_k_index[13559] = 63338;
mem_k_index[13560] = 63341;
mem_k_index[13561] = 63343;
mem_k_index[13562] = 63346;
mem_k_index[13563] = 63348;
mem_k_index[13564] = 63351;
mem_k_index[13565] = 63353;
mem_k_index[13566] = 63356;
mem_k_index[13567] = 63358;
mem_k_index[13568] = 63680;
mem_k_index[13569] = 63682;
mem_k_index[13570] = 63685;
mem_k_index[13571] = 63687;
mem_k_index[13572] = 63690;
mem_k_index[13573] = 63692;
mem_k_index[13574] = 63695;
mem_k_index[13575] = 63697;
mem_k_index[13576] = 63700;
mem_k_index[13577] = 63702;
mem_k_index[13578] = 63705;
mem_k_index[13579] = 63707;
mem_k_index[13580] = 63710;
mem_k_index[13581] = 63712;
mem_k_index[13582] = 63715;
mem_k_index[13583] = 63717;
mem_k_index[13584] = 63720;
mem_k_index[13585] = 63722;
mem_k_index[13586] = 63725;
mem_k_index[13587] = 63727;
mem_k_index[13588] = 63730;
mem_k_index[13589] = 63732;
mem_k_index[13590] = 63735;
mem_k_index[13591] = 63737;
mem_k_index[13592] = 63740;
mem_k_index[13593] = 63742;
mem_k_index[13594] = 63745;
mem_k_index[13595] = 63747;
mem_k_index[13596] = 63750;
mem_k_index[13597] = 63752;
mem_k_index[13598] = 63755;
mem_k_index[13599] = 63757;
mem_k_index[13600] = 63760;
mem_k_index[13601] = 63762;
mem_k_index[13602] = 63765;
mem_k_index[13603] = 63767;
mem_k_index[13604] = 63770;
mem_k_index[13605] = 63772;
mem_k_index[13606] = 63775;
mem_k_index[13607] = 63777;
mem_k_index[13608] = 63780;
mem_k_index[13609] = 63782;
mem_k_index[13610] = 63785;
mem_k_index[13611] = 63788;
mem_k_index[13612] = 63790;
mem_k_index[13613] = 63793;
mem_k_index[13614] = 63795;
mem_k_index[13615] = 63798;
mem_k_index[13616] = 63800;
mem_k_index[13617] = 63803;
mem_k_index[13618] = 63805;
mem_k_index[13619] = 63808;
mem_k_index[13620] = 63810;
mem_k_index[13621] = 63813;
mem_k_index[13622] = 63815;
mem_k_index[13623] = 63818;
mem_k_index[13624] = 63820;
mem_k_index[13625] = 63823;
mem_k_index[13626] = 63825;
mem_k_index[13627] = 63828;
mem_k_index[13628] = 63830;
mem_k_index[13629] = 63833;
mem_k_index[13630] = 63835;
mem_k_index[13631] = 63838;
mem_k_index[13632] = 63840;
mem_k_index[13633] = 63843;
mem_k_index[13634] = 63845;
mem_k_index[13635] = 63848;
mem_k_index[13636] = 63850;
mem_k_index[13637] = 63853;
mem_k_index[13638] = 63855;
mem_k_index[13639] = 63858;
mem_k_index[13640] = 63860;
mem_k_index[13641] = 63863;
mem_k_index[13642] = 63865;
mem_k_index[13643] = 63868;
mem_k_index[13644] = 63870;
mem_k_index[13645] = 63873;
mem_k_index[13646] = 63875;
mem_k_index[13647] = 63878;
mem_k_index[13648] = 63880;
mem_k_index[13649] = 63883;
mem_k_index[13650] = 63885;
mem_k_index[13651] = 63888;
mem_k_index[13652] = 63890;
mem_k_index[13653] = 63893;
mem_k_index[13654] = 63896;
mem_k_index[13655] = 63898;
mem_k_index[13656] = 63901;
mem_k_index[13657] = 63903;
mem_k_index[13658] = 63906;
mem_k_index[13659] = 63908;
mem_k_index[13660] = 63911;
mem_k_index[13661] = 63913;
mem_k_index[13662] = 63916;
mem_k_index[13663] = 63918;
mem_k_index[13664] = 63921;
mem_k_index[13665] = 63923;
mem_k_index[13666] = 63926;
mem_k_index[13667] = 63928;
mem_k_index[13668] = 63931;
mem_k_index[13669] = 63933;
mem_k_index[13670] = 63936;
mem_k_index[13671] = 63938;
mem_k_index[13672] = 63941;
mem_k_index[13673] = 63943;
mem_k_index[13674] = 63946;
mem_k_index[13675] = 63948;
mem_k_index[13676] = 63951;
mem_k_index[13677] = 63953;
mem_k_index[13678] = 63956;
mem_k_index[13679] = 63958;
mem_k_index[13680] = 63961;
mem_k_index[13681] = 63963;
mem_k_index[13682] = 63966;
mem_k_index[13683] = 63968;
mem_k_index[13684] = 63971;
mem_k_index[13685] = 63973;
mem_k_index[13686] = 63976;
mem_k_index[13687] = 63978;
mem_k_index[13688] = 63981;
mem_k_index[13689] = 63983;
mem_k_index[13690] = 63986;
mem_k_index[13691] = 63988;
mem_k_index[13692] = 63991;
mem_k_index[13693] = 63993;
mem_k_index[13694] = 63996;
mem_k_index[13695] = 63998;
mem_k_index[13696] = 64320;
mem_k_index[13697] = 64322;
mem_k_index[13698] = 64325;
mem_k_index[13699] = 64327;
mem_k_index[13700] = 64330;
mem_k_index[13701] = 64332;
mem_k_index[13702] = 64335;
mem_k_index[13703] = 64337;
mem_k_index[13704] = 64340;
mem_k_index[13705] = 64342;
mem_k_index[13706] = 64345;
mem_k_index[13707] = 64347;
mem_k_index[13708] = 64350;
mem_k_index[13709] = 64352;
mem_k_index[13710] = 64355;
mem_k_index[13711] = 64357;
mem_k_index[13712] = 64360;
mem_k_index[13713] = 64362;
mem_k_index[13714] = 64365;
mem_k_index[13715] = 64367;
mem_k_index[13716] = 64370;
mem_k_index[13717] = 64372;
mem_k_index[13718] = 64375;
mem_k_index[13719] = 64377;
mem_k_index[13720] = 64380;
mem_k_index[13721] = 64382;
mem_k_index[13722] = 64385;
mem_k_index[13723] = 64387;
mem_k_index[13724] = 64390;
mem_k_index[13725] = 64392;
mem_k_index[13726] = 64395;
mem_k_index[13727] = 64397;
mem_k_index[13728] = 64400;
mem_k_index[13729] = 64402;
mem_k_index[13730] = 64405;
mem_k_index[13731] = 64407;
mem_k_index[13732] = 64410;
mem_k_index[13733] = 64412;
mem_k_index[13734] = 64415;
mem_k_index[13735] = 64417;
mem_k_index[13736] = 64420;
mem_k_index[13737] = 64422;
mem_k_index[13738] = 64425;
mem_k_index[13739] = 64428;
mem_k_index[13740] = 64430;
mem_k_index[13741] = 64433;
mem_k_index[13742] = 64435;
mem_k_index[13743] = 64438;
mem_k_index[13744] = 64440;
mem_k_index[13745] = 64443;
mem_k_index[13746] = 64445;
mem_k_index[13747] = 64448;
mem_k_index[13748] = 64450;
mem_k_index[13749] = 64453;
mem_k_index[13750] = 64455;
mem_k_index[13751] = 64458;
mem_k_index[13752] = 64460;
mem_k_index[13753] = 64463;
mem_k_index[13754] = 64465;
mem_k_index[13755] = 64468;
mem_k_index[13756] = 64470;
mem_k_index[13757] = 64473;
mem_k_index[13758] = 64475;
mem_k_index[13759] = 64478;
mem_k_index[13760] = 64480;
mem_k_index[13761] = 64483;
mem_k_index[13762] = 64485;
mem_k_index[13763] = 64488;
mem_k_index[13764] = 64490;
mem_k_index[13765] = 64493;
mem_k_index[13766] = 64495;
mem_k_index[13767] = 64498;
mem_k_index[13768] = 64500;
mem_k_index[13769] = 64503;
mem_k_index[13770] = 64505;
mem_k_index[13771] = 64508;
mem_k_index[13772] = 64510;
mem_k_index[13773] = 64513;
mem_k_index[13774] = 64515;
mem_k_index[13775] = 64518;
mem_k_index[13776] = 64520;
mem_k_index[13777] = 64523;
mem_k_index[13778] = 64525;
mem_k_index[13779] = 64528;
mem_k_index[13780] = 64530;
mem_k_index[13781] = 64533;
mem_k_index[13782] = 64536;
mem_k_index[13783] = 64538;
mem_k_index[13784] = 64541;
mem_k_index[13785] = 64543;
mem_k_index[13786] = 64546;
mem_k_index[13787] = 64548;
mem_k_index[13788] = 64551;
mem_k_index[13789] = 64553;
mem_k_index[13790] = 64556;
mem_k_index[13791] = 64558;
mem_k_index[13792] = 64561;
mem_k_index[13793] = 64563;
mem_k_index[13794] = 64566;
mem_k_index[13795] = 64568;
mem_k_index[13796] = 64571;
mem_k_index[13797] = 64573;
mem_k_index[13798] = 64576;
mem_k_index[13799] = 64578;
mem_k_index[13800] = 64581;
mem_k_index[13801] = 64583;
mem_k_index[13802] = 64586;
mem_k_index[13803] = 64588;
mem_k_index[13804] = 64591;
mem_k_index[13805] = 64593;
mem_k_index[13806] = 64596;
mem_k_index[13807] = 64598;
mem_k_index[13808] = 64601;
mem_k_index[13809] = 64603;
mem_k_index[13810] = 64606;
mem_k_index[13811] = 64608;
mem_k_index[13812] = 64611;
mem_k_index[13813] = 64613;
mem_k_index[13814] = 64616;
mem_k_index[13815] = 64618;
mem_k_index[13816] = 64621;
mem_k_index[13817] = 64623;
mem_k_index[13818] = 64626;
mem_k_index[13819] = 64628;
mem_k_index[13820] = 64631;
mem_k_index[13821] = 64633;
mem_k_index[13822] = 64636;
mem_k_index[13823] = 64638;
mem_k_index[13824] = 64960;
mem_k_index[13825] = 64962;
mem_k_index[13826] = 64965;
mem_k_index[13827] = 64967;
mem_k_index[13828] = 64970;
mem_k_index[13829] = 64972;
mem_k_index[13830] = 64975;
mem_k_index[13831] = 64977;
mem_k_index[13832] = 64980;
mem_k_index[13833] = 64982;
mem_k_index[13834] = 64985;
mem_k_index[13835] = 64987;
mem_k_index[13836] = 64990;
mem_k_index[13837] = 64992;
mem_k_index[13838] = 64995;
mem_k_index[13839] = 64997;
mem_k_index[13840] = 65000;
mem_k_index[13841] = 65002;
mem_k_index[13842] = 65005;
mem_k_index[13843] = 65007;
mem_k_index[13844] = 65010;
mem_k_index[13845] = 65012;
mem_k_index[13846] = 65015;
mem_k_index[13847] = 65017;
mem_k_index[13848] = 65020;
mem_k_index[13849] = 65022;
mem_k_index[13850] = 65025;
mem_k_index[13851] = 65027;
mem_k_index[13852] = 65030;
mem_k_index[13853] = 65032;
mem_k_index[13854] = 65035;
mem_k_index[13855] = 65037;
mem_k_index[13856] = 65040;
mem_k_index[13857] = 65042;
mem_k_index[13858] = 65045;
mem_k_index[13859] = 65047;
mem_k_index[13860] = 65050;
mem_k_index[13861] = 65052;
mem_k_index[13862] = 65055;
mem_k_index[13863] = 65057;
mem_k_index[13864] = 65060;
mem_k_index[13865] = 65062;
mem_k_index[13866] = 65065;
mem_k_index[13867] = 65068;
mem_k_index[13868] = 65070;
mem_k_index[13869] = 65073;
mem_k_index[13870] = 65075;
mem_k_index[13871] = 65078;
mem_k_index[13872] = 65080;
mem_k_index[13873] = 65083;
mem_k_index[13874] = 65085;
mem_k_index[13875] = 65088;
mem_k_index[13876] = 65090;
mem_k_index[13877] = 65093;
mem_k_index[13878] = 65095;
mem_k_index[13879] = 65098;
mem_k_index[13880] = 65100;
mem_k_index[13881] = 65103;
mem_k_index[13882] = 65105;
mem_k_index[13883] = 65108;
mem_k_index[13884] = 65110;
mem_k_index[13885] = 65113;
mem_k_index[13886] = 65115;
mem_k_index[13887] = 65118;
mem_k_index[13888] = 65120;
mem_k_index[13889] = 65123;
mem_k_index[13890] = 65125;
mem_k_index[13891] = 65128;
mem_k_index[13892] = 65130;
mem_k_index[13893] = 65133;
mem_k_index[13894] = 65135;
mem_k_index[13895] = 65138;
mem_k_index[13896] = 65140;
mem_k_index[13897] = 65143;
mem_k_index[13898] = 65145;
mem_k_index[13899] = 65148;
mem_k_index[13900] = 65150;
mem_k_index[13901] = 65153;
mem_k_index[13902] = 65155;
mem_k_index[13903] = 65158;
mem_k_index[13904] = 65160;
mem_k_index[13905] = 65163;
mem_k_index[13906] = 65165;
mem_k_index[13907] = 65168;
mem_k_index[13908] = 65170;
mem_k_index[13909] = 65173;
mem_k_index[13910] = 65176;
mem_k_index[13911] = 65178;
mem_k_index[13912] = 65181;
mem_k_index[13913] = 65183;
mem_k_index[13914] = 65186;
mem_k_index[13915] = 65188;
mem_k_index[13916] = 65191;
mem_k_index[13917] = 65193;
mem_k_index[13918] = 65196;
mem_k_index[13919] = 65198;
mem_k_index[13920] = 65201;
mem_k_index[13921] = 65203;
mem_k_index[13922] = 65206;
mem_k_index[13923] = 65208;
mem_k_index[13924] = 65211;
mem_k_index[13925] = 65213;
mem_k_index[13926] = 65216;
mem_k_index[13927] = 65218;
mem_k_index[13928] = 65221;
mem_k_index[13929] = 65223;
mem_k_index[13930] = 65226;
mem_k_index[13931] = 65228;
mem_k_index[13932] = 65231;
mem_k_index[13933] = 65233;
mem_k_index[13934] = 65236;
mem_k_index[13935] = 65238;
mem_k_index[13936] = 65241;
mem_k_index[13937] = 65243;
mem_k_index[13938] = 65246;
mem_k_index[13939] = 65248;
mem_k_index[13940] = 65251;
mem_k_index[13941] = 65253;
mem_k_index[13942] = 65256;
mem_k_index[13943] = 65258;
mem_k_index[13944] = 65261;
mem_k_index[13945] = 65263;
mem_k_index[13946] = 65266;
mem_k_index[13947] = 65268;
mem_k_index[13948] = 65271;
mem_k_index[13949] = 65273;
mem_k_index[13950] = 65276;
mem_k_index[13951] = 65278;
mem_k_index[13952] = 65600;
mem_k_index[13953] = 65602;
mem_k_index[13954] = 65605;
mem_k_index[13955] = 65607;
mem_k_index[13956] = 65610;
mem_k_index[13957] = 65612;
mem_k_index[13958] = 65615;
mem_k_index[13959] = 65617;
mem_k_index[13960] = 65620;
mem_k_index[13961] = 65622;
mem_k_index[13962] = 65625;
mem_k_index[13963] = 65627;
mem_k_index[13964] = 65630;
mem_k_index[13965] = 65632;
mem_k_index[13966] = 65635;
mem_k_index[13967] = 65637;
mem_k_index[13968] = 65640;
mem_k_index[13969] = 65642;
mem_k_index[13970] = 65645;
mem_k_index[13971] = 65647;
mem_k_index[13972] = 65650;
mem_k_index[13973] = 65652;
mem_k_index[13974] = 65655;
mem_k_index[13975] = 65657;
mem_k_index[13976] = 65660;
mem_k_index[13977] = 65662;
mem_k_index[13978] = 65665;
mem_k_index[13979] = 65667;
mem_k_index[13980] = 65670;
mem_k_index[13981] = 65672;
mem_k_index[13982] = 65675;
mem_k_index[13983] = 65677;
mem_k_index[13984] = 65680;
mem_k_index[13985] = 65682;
mem_k_index[13986] = 65685;
mem_k_index[13987] = 65687;
mem_k_index[13988] = 65690;
mem_k_index[13989] = 65692;
mem_k_index[13990] = 65695;
mem_k_index[13991] = 65697;
mem_k_index[13992] = 65700;
mem_k_index[13993] = 65702;
mem_k_index[13994] = 65705;
mem_k_index[13995] = 65708;
mem_k_index[13996] = 65710;
mem_k_index[13997] = 65713;
mem_k_index[13998] = 65715;
mem_k_index[13999] = 65718;
mem_k_index[14000] = 65720;
mem_k_index[14001] = 65723;
mem_k_index[14002] = 65725;
mem_k_index[14003] = 65728;
mem_k_index[14004] = 65730;
mem_k_index[14005] = 65733;
mem_k_index[14006] = 65735;
mem_k_index[14007] = 65738;
mem_k_index[14008] = 65740;
mem_k_index[14009] = 65743;
mem_k_index[14010] = 65745;
mem_k_index[14011] = 65748;
mem_k_index[14012] = 65750;
mem_k_index[14013] = 65753;
mem_k_index[14014] = 65755;
mem_k_index[14015] = 65758;
mem_k_index[14016] = 65760;
mem_k_index[14017] = 65763;
mem_k_index[14018] = 65765;
mem_k_index[14019] = 65768;
mem_k_index[14020] = 65770;
mem_k_index[14021] = 65773;
mem_k_index[14022] = 65775;
mem_k_index[14023] = 65778;
mem_k_index[14024] = 65780;
mem_k_index[14025] = 65783;
mem_k_index[14026] = 65785;
mem_k_index[14027] = 65788;
mem_k_index[14028] = 65790;
mem_k_index[14029] = 65793;
mem_k_index[14030] = 65795;
mem_k_index[14031] = 65798;
mem_k_index[14032] = 65800;
mem_k_index[14033] = 65803;
mem_k_index[14034] = 65805;
mem_k_index[14035] = 65808;
mem_k_index[14036] = 65810;
mem_k_index[14037] = 65813;
mem_k_index[14038] = 65816;
mem_k_index[14039] = 65818;
mem_k_index[14040] = 65821;
mem_k_index[14041] = 65823;
mem_k_index[14042] = 65826;
mem_k_index[14043] = 65828;
mem_k_index[14044] = 65831;
mem_k_index[14045] = 65833;
mem_k_index[14046] = 65836;
mem_k_index[14047] = 65838;
mem_k_index[14048] = 65841;
mem_k_index[14049] = 65843;
mem_k_index[14050] = 65846;
mem_k_index[14051] = 65848;
mem_k_index[14052] = 65851;
mem_k_index[14053] = 65853;
mem_k_index[14054] = 65856;
mem_k_index[14055] = 65858;
mem_k_index[14056] = 65861;
mem_k_index[14057] = 65863;
mem_k_index[14058] = 65866;
mem_k_index[14059] = 65868;
mem_k_index[14060] = 65871;
mem_k_index[14061] = 65873;
mem_k_index[14062] = 65876;
mem_k_index[14063] = 65878;
mem_k_index[14064] = 65881;
mem_k_index[14065] = 65883;
mem_k_index[14066] = 65886;
mem_k_index[14067] = 65888;
mem_k_index[14068] = 65891;
mem_k_index[14069] = 65893;
mem_k_index[14070] = 65896;
mem_k_index[14071] = 65898;
mem_k_index[14072] = 65901;
mem_k_index[14073] = 65903;
mem_k_index[14074] = 65906;
mem_k_index[14075] = 65908;
mem_k_index[14076] = 65911;
mem_k_index[14077] = 65913;
mem_k_index[14078] = 65916;
mem_k_index[14079] = 65918;
mem_k_index[14080] = 66240;
mem_k_index[14081] = 66242;
mem_k_index[14082] = 66245;
mem_k_index[14083] = 66247;
mem_k_index[14084] = 66250;
mem_k_index[14085] = 66252;
mem_k_index[14086] = 66255;
mem_k_index[14087] = 66257;
mem_k_index[14088] = 66260;
mem_k_index[14089] = 66262;
mem_k_index[14090] = 66265;
mem_k_index[14091] = 66267;
mem_k_index[14092] = 66270;
mem_k_index[14093] = 66272;
mem_k_index[14094] = 66275;
mem_k_index[14095] = 66277;
mem_k_index[14096] = 66280;
mem_k_index[14097] = 66282;
mem_k_index[14098] = 66285;
mem_k_index[14099] = 66287;
mem_k_index[14100] = 66290;
mem_k_index[14101] = 66292;
mem_k_index[14102] = 66295;
mem_k_index[14103] = 66297;
mem_k_index[14104] = 66300;
mem_k_index[14105] = 66302;
mem_k_index[14106] = 66305;
mem_k_index[14107] = 66307;
mem_k_index[14108] = 66310;
mem_k_index[14109] = 66312;
mem_k_index[14110] = 66315;
mem_k_index[14111] = 66317;
mem_k_index[14112] = 66320;
mem_k_index[14113] = 66322;
mem_k_index[14114] = 66325;
mem_k_index[14115] = 66327;
mem_k_index[14116] = 66330;
mem_k_index[14117] = 66332;
mem_k_index[14118] = 66335;
mem_k_index[14119] = 66337;
mem_k_index[14120] = 66340;
mem_k_index[14121] = 66342;
mem_k_index[14122] = 66345;
mem_k_index[14123] = 66348;
mem_k_index[14124] = 66350;
mem_k_index[14125] = 66353;
mem_k_index[14126] = 66355;
mem_k_index[14127] = 66358;
mem_k_index[14128] = 66360;
mem_k_index[14129] = 66363;
mem_k_index[14130] = 66365;
mem_k_index[14131] = 66368;
mem_k_index[14132] = 66370;
mem_k_index[14133] = 66373;
mem_k_index[14134] = 66375;
mem_k_index[14135] = 66378;
mem_k_index[14136] = 66380;
mem_k_index[14137] = 66383;
mem_k_index[14138] = 66385;
mem_k_index[14139] = 66388;
mem_k_index[14140] = 66390;
mem_k_index[14141] = 66393;
mem_k_index[14142] = 66395;
mem_k_index[14143] = 66398;
mem_k_index[14144] = 66400;
mem_k_index[14145] = 66403;
mem_k_index[14146] = 66405;
mem_k_index[14147] = 66408;
mem_k_index[14148] = 66410;
mem_k_index[14149] = 66413;
mem_k_index[14150] = 66415;
mem_k_index[14151] = 66418;
mem_k_index[14152] = 66420;
mem_k_index[14153] = 66423;
mem_k_index[14154] = 66425;
mem_k_index[14155] = 66428;
mem_k_index[14156] = 66430;
mem_k_index[14157] = 66433;
mem_k_index[14158] = 66435;
mem_k_index[14159] = 66438;
mem_k_index[14160] = 66440;
mem_k_index[14161] = 66443;
mem_k_index[14162] = 66445;
mem_k_index[14163] = 66448;
mem_k_index[14164] = 66450;
mem_k_index[14165] = 66453;
mem_k_index[14166] = 66456;
mem_k_index[14167] = 66458;
mem_k_index[14168] = 66461;
mem_k_index[14169] = 66463;
mem_k_index[14170] = 66466;
mem_k_index[14171] = 66468;
mem_k_index[14172] = 66471;
mem_k_index[14173] = 66473;
mem_k_index[14174] = 66476;
mem_k_index[14175] = 66478;
mem_k_index[14176] = 66481;
mem_k_index[14177] = 66483;
mem_k_index[14178] = 66486;
mem_k_index[14179] = 66488;
mem_k_index[14180] = 66491;
mem_k_index[14181] = 66493;
mem_k_index[14182] = 66496;
mem_k_index[14183] = 66498;
mem_k_index[14184] = 66501;
mem_k_index[14185] = 66503;
mem_k_index[14186] = 66506;
mem_k_index[14187] = 66508;
mem_k_index[14188] = 66511;
mem_k_index[14189] = 66513;
mem_k_index[14190] = 66516;
mem_k_index[14191] = 66518;
mem_k_index[14192] = 66521;
mem_k_index[14193] = 66523;
mem_k_index[14194] = 66526;
mem_k_index[14195] = 66528;
mem_k_index[14196] = 66531;
mem_k_index[14197] = 66533;
mem_k_index[14198] = 66536;
mem_k_index[14199] = 66538;
mem_k_index[14200] = 66541;
mem_k_index[14201] = 66543;
mem_k_index[14202] = 66546;
mem_k_index[14203] = 66548;
mem_k_index[14204] = 66551;
mem_k_index[14205] = 66553;
mem_k_index[14206] = 66556;
mem_k_index[14207] = 66558;
mem_k_index[14208] = 66560;
mem_k_index[14209] = 66562;
mem_k_index[14210] = 66565;
mem_k_index[14211] = 66567;
mem_k_index[14212] = 66570;
mem_k_index[14213] = 66572;
mem_k_index[14214] = 66575;
mem_k_index[14215] = 66577;
mem_k_index[14216] = 66580;
mem_k_index[14217] = 66582;
mem_k_index[14218] = 66585;
mem_k_index[14219] = 66587;
mem_k_index[14220] = 66590;
mem_k_index[14221] = 66592;
mem_k_index[14222] = 66595;
mem_k_index[14223] = 66597;
mem_k_index[14224] = 66600;
mem_k_index[14225] = 66602;
mem_k_index[14226] = 66605;
mem_k_index[14227] = 66607;
mem_k_index[14228] = 66610;
mem_k_index[14229] = 66612;
mem_k_index[14230] = 66615;
mem_k_index[14231] = 66617;
mem_k_index[14232] = 66620;
mem_k_index[14233] = 66622;
mem_k_index[14234] = 66625;
mem_k_index[14235] = 66627;
mem_k_index[14236] = 66630;
mem_k_index[14237] = 66632;
mem_k_index[14238] = 66635;
mem_k_index[14239] = 66637;
mem_k_index[14240] = 66640;
mem_k_index[14241] = 66642;
mem_k_index[14242] = 66645;
mem_k_index[14243] = 66647;
mem_k_index[14244] = 66650;
mem_k_index[14245] = 66652;
mem_k_index[14246] = 66655;
mem_k_index[14247] = 66657;
mem_k_index[14248] = 66660;
mem_k_index[14249] = 66662;
mem_k_index[14250] = 66665;
mem_k_index[14251] = 66668;
mem_k_index[14252] = 66670;
mem_k_index[14253] = 66673;
mem_k_index[14254] = 66675;
mem_k_index[14255] = 66678;
mem_k_index[14256] = 66680;
mem_k_index[14257] = 66683;
mem_k_index[14258] = 66685;
mem_k_index[14259] = 66688;
mem_k_index[14260] = 66690;
mem_k_index[14261] = 66693;
mem_k_index[14262] = 66695;
mem_k_index[14263] = 66698;
mem_k_index[14264] = 66700;
mem_k_index[14265] = 66703;
mem_k_index[14266] = 66705;
mem_k_index[14267] = 66708;
mem_k_index[14268] = 66710;
mem_k_index[14269] = 66713;
mem_k_index[14270] = 66715;
mem_k_index[14271] = 66718;
mem_k_index[14272] = 66720;
mem_k_index[14273] = 66723;
mem_k_index[14274] = 66725;
mem_k_index[14275] = 66728;
mem_k_index[14276] = 66730;
mem_k_index[14277] = 66733;
mem_k_index[14278] = 66735;
mem_k_index[14279] = 66738;
mem_k_index[14280] = 66740;
mem_k_index[14281] = 66743;
mem_k_index[14282] = 66745;
mem_k_index[14283] = 66748;
mem_k_index[14284] = 66750;
mem_k_index[14285] = 66753;
mem_k_index[14286] = 66755;
mem_k_index[14287] = 66758;
mem_k_index[14288] = 66760;
mem_k_index[14289] = 66763;
mem_k_index[14290] = 66765;
mem_k_index[14291] = 66768;
mem_k_index[14292] = 66770;
mem_k_index[14293] = 66773;
mem_k_index[14294] = 66776;
mem_k_index[14295] = 66778;
mem_k_index[14296] = 66781;
mem_k_index[14297] = 66783;
mem_k_index[14298] = 66786;
mem_k_index[14299] = 66788;
mem_k_index[14300] = 66791;
mem_k_index[14301] = 66793;
mem_k_index[14302] = 66796;
mem_k_index[14303] = 66798;
mem_k_index[14304] = 66801;
mem_k_index[14305] = 66803;
mem_k_index[14306] = 66806;
mem_k_index[14307] = 66808;
mem_k_index[14308] = 66811;
mem_k_index[14309] = 66813;
mem_k_index[14310] = 66816;
mem_k_index[14311] = 66818;
mem_k_index[14312] = 66821;
mem_k_index[14313] = 66823;
mem_k_index[14314] = 66826;
mem_k_index[14315] = 66828;
mem_k_index[14316] = 66831;
mem_k_index[14317] = 66833;
mem_k_index[14318] = 66836;
mem_k_index[14319] = 66838;
mem_k_index[14320] = 66841;
mem_k_index[14321] = 66843;
mem_k_index[14322] = 66846;
mem_k_index[14323] = 66848;
mem_k_index[14324] = 66851;
mem_k_index[14325] = 66853;
mem_k_index[14326] = 66856;
mem_k_index[14327] = 66858;
mem_k_index[14328] = 66861;
mem_k_index[14329] = 66863;
mem_k_index[14330] = 66866;
mem_k_index[14331] = 66868;
mem_k_index[14332] = 66871;
mem_k_index[14333] = 66873;
mem_k_index[14334] = 66876;
mem_k_index[14335] = 66878;
mem_k_index[14336] = 67200;
mem_k_index[14337] = 67202;
mem_k_index[14338] = 67205;
mem_k_index[14339] = 67207;
mem_k_index[14340] = 67210;
mem_k_index[14341] = 67212;
mem_k_index[14342] = 67215;
mem_k_index[14343] = 67217;
mem_k_index[14344] = 67220;
mem_k_index[14345] = 67222;
mem_k_index[14346] = 67225;
mem_k_index[14347] = 67227;
mem_k_index[14348] = 67230;
mem_k_index[14349] = 67232;
mem_k_index[14350] = 67235;
mem_k_index[14351] = 67237;
mem_k_index[14352] = 67240;
mem_k_index[14353] = 67242;
mem_k_index[14354] = 67245;
mem_k_index[14355] = 67247;
mem_k_index[14356] = 67250;
mem_k_index[14357] = 67252;
mem_k_index[14358] = 67255;
mem_k_index[14359] = 67257;
mem_k_index[14360] = 67260;
mem_k_index[14361] = 67262;
mem_k_index[14362] = 67265;
mem_k_index[14363] = 67267;
mem_k_index[14364] = 67270;
mem_k_index[14365] = 67272;
mem_k_index[14366] = 67275;
mem_k_index[14367] = 67277;
mem_k_index[14368] = 67280;
mem_k_index[14369] = 67282;
mem_k_index[14370] = 67285;
mem_k_index[14371] = 67287;
mem_k_index[14372] = 67290;
mem_k_index[14373] = 67292;
mem_k_index[14374] = 67295;
mem_k_index[14375] = 67297;
mem_k_index[14376] = 67300;
mem_k_index[14377] = 67302;
mem_k_index[14378] = 67305;
mem_k_index[14379] = 67308;
mem_k_index[14380] = 67310;
mem_k_index[14381] = 67313;
mem_k_index[14382] = 67315;
mem_k_index[14383] = 67318;
mem_k_index[14384] = 67320;
mem_k_index[14385] = 67323;
mem_k_index[14386] = 67325;
mem_k_index[14387] = 67328;
mem_k_index[14388] = 67330;
mem_k_index[14389] = 67333;
mem_k_index[14390] = 67335;
mem_k_index[14391] = 67338;
mem_k_index[14392] = 67340;
mem_k_index[14393] = 67343;
mem_k_index[14394] = 67345;
mem_k_index[14395] = 67348;
mem_k_index[14396] = 67350;
mem_k_index[14397] = 67353;
mem_k_index[14398] = 67355;
mem_k_index[14399] = 67358;
mem_k_index[14400] = 67360;
mem_k_index[14401] = 67363;
mem_k_index[14402] = 67365;
mem_k_index[14403] = 67368;
mem_k_index[14404] = 67370;
mem_k_index[14405] = 67373;
mem_k_index[14406] = 67375;
mem_k_index[14407] = 67378;
mem_k_index[14408] = 67380;
mem_k_index[14409] = 67383;
mem_k_index[14410] = 67385;
mem_k_index[14411] = 67388;
mem_k_index[14412] = 67390;
mem_k_index[14413] = 67393;
mem_k_index[14414] = 67395;
mem_k_index[14415] = 67398;
mem_k_index[14416] = 67400;
mem_k_index[14417] = 67403;
mem_k_index[14418] = 67405;
mem_k_index[14419] = 67408;
mem_k_index[14420] = 67410;
mem_k_index[14421] = 67413;
mem_k_index[14422] = 67416;
mem_k_index[14423] = 67418;
mem_k_index[14424] = 67421;
mem_k_index[14425] = 67423;
mem_k_index[14426] = 67426;
mem_k_index[14427] = 67428;
mem_k_index[14428] = 67431;
mem_k_index[14429] = 67433;
mem_k_index[14430] = 67436;
mem_k_index[14431] = 67438;
mem_k_index[14432] = 67441;
mem_k_index[14433] = 67443;
mem_k_index[14434] = 67446;
mem_k_index[14435] = 67448;
mem_k_index[14436] = 67451;
mem_k_index[14437] = 67453;
mem_k_index[14438] = 67456;
mem_k_index[14439] = 67458;
mem_k_index[14440] = 67461;
mem_k_index[14441] = 67463;
mem_k_index[14442] = 67466;
mem_k_index[14443] = 67468;
mem_k_index[14444] = 67471;
mem_k_index[14445] = 67473;
mem_k_index[14446] = 67476;
mem_k_index[14447] = 67478;
mem_k_index[14448] = 67481;
mem_k_index[14449] = 67483;
mem_k_index[14450] = 67486;
mem_k_index[14451] = 67488;
mem_k_index[14452] = 67491;
mem_k_index[14453] = 67493;
mem_k_index[14454] = 67496;
mem_k_index[14455] = 67498;
mem_k_index[14456] = 67501;
mem_k_index[14457] = 67503;
mem_k_index[14458] = 67506;
mem_k_index[14459] = 67508;
mem_k_index[14460] = 67511;
mem_k_index[14461] = 67513;
mem_k_index[14462] = 67516;
mem_k_index[14463] = 67518;
mem_k_index[14464] = 67840;
mem_k_index[14465] = 67842;
mem_k_index[14466] = 67845;
mem_k_index[14467] = 67847;
mem_k_index[14468] = 67850;
mem_k_index[14469] = 67852;
mem_k_index[14470] = 67855;
mem_k_index[14471] = 67857;
mem_k_index[14472] = 67860;
mem_k_index[14473] = 67862;
mem_k_index[14474] = 67865;
mem_k_index[14475] = 67867;
mem_k_index[14476] = 67870;
mem_k_index[14477] = 67872;
mem_k_index[14478] = 67875;
mem_k_index[14479] = 67877;
mem_k_index[14480] = 67880;
mem_k_index[14481] = 67882;
mem_k_index[14482] = 67885;
mem_k_index[14483] = 67887;
mem_k_index[14484] = 67890;
mem_k_index[14485] = 67892;
mem_k_index[14486] = 67895;
mem_k_index[14487] = 67897;
mem_k_index[14488] = 67900;
mem_k_index[14489] = 67902;
mem_k_index[14490] = 67905;
mem_k_index[14491] = 67907;
mem_k_index[14492] = 67910;
mem_k_index[14493] = 67912;
mem_k_index[14494] = 67915;
mem_k_index[14495] = 67917;
mem_k_index[14496] = 67920;
mem_k_index[14497] = 67922;
mem_k_index[14498] = 67925;
mem_k_index[14499] = 67927;
mem_k_index[14500] = 67930;
mem_k_index[14501] = 67932;
mem_k_index[14502] = 67935;
mem_k_index[14503] = 67937;
mem_k_index[14504] = 67940;
mem_k_index[14505] = 67942;
mem_k_index[14506] = 67945;
mem_k_index[14507] = 67948;
mem_k_index[14508] = 67950;
mem_k_index[14509] = 67953;
mem_k_index[14510] = 67955;
mem_k_index[14511] = 67958;
mem_k_index[14512] = 67960;
mem_k_index[14513] = 67963;
mem_k_index[14514] = 67965;
mem_k_index[14515] = 67968;
mem_k_index[14516] = 67970;
mem_k_index[14517] = 67973;
mem_k_index[14518] = 67975;
mem_k_index[14519] = 67978;
mem_k_index[14520] = 67980;
mem_k_index[14521] = 67983;
mem_k_index[14522] = 67985;
mem_k_index[14523] = 67988;
mem_k_index[14524] = 67990;
mem_k_index[14525] = 67993;
mem_k_index[14526] = 67995;
mem_k_index[14527] = 67998;
mem_k_index[14528] = 68000;
mem_k_index[14529] = 68003;
mem_k_index[14530] = 68005;
mem_k_index[14531] = 68008;
mem_k_index[14532] = 68010;
mem_k_index[14533] = 68013;
mem_k_index[14534] = 68015;
mem_k_index[14535] = 68018;
mem_k_index[14536] = 68020;
mem_k_index[14537] = 68023;
mem_k_index[14538] = 68025;
mem_k_index[14539] = 68028;
mem_k_index[14540] = 68030;
mem_k_index[14541] = 68033;
mem_k_index[14542] = 68035;
mem_k_index[14543] = 68038;
mem_k_index[14544] = 68040;
mem_k_index[14545] = 68043;
mem_k_index[14546] = 68045;
mem_k_index[14547] = 68048;
mem_k_index[14548] = 68050;
mem_k_index[14549] = 68053;
mem_k_index[14550] = 68056;
mem_k_index[14551] = 68058;
mem_k_index[14552] = 68061;
mem_k_index[14553] = 68063;
mem_k_index[14554] = 68066;
mem_k_index[14555] = 68068;
mem_k_index[14556] = 68071;
mem_k_index[14557] = 68073;
mem_k_index[14558] = 68076;
mem_k_index[14559] = 68078;
mem_k_index[14560] = 68081;
mem_k_index[14561] = 68083;
mem_k_index[14562] = 68086;
mem_k_index[14563] = 68088;
mem_k_index[14564] = 68091;
mem_k_index[14565] = 68093;
mem_k_index[14566] = 68096;
mem_k_index[14567] = 68098;
mem_k_index[14568] = 68101;
mem_k_index[14569] = 68103;
mem_k_index[14570] = 68106;
mem_k_index[14571] = 68108;
mem_k_index[14572] = 68111;
mem_k_index[14573] = 68113;
mem_k_index[14574] = 68116;
mem_k_index[14575] = 68118;
mem_k_index[14576] = 68121;
mem_k_index[14577] = 68123;
mem_k_index[14578] = 68126;
mem_k_index[14579] = 68128;
mem_k_index[14580] = 68131;
mem_k_index[14581] = 68133;
mem_k_index[14582] = 68136;
mem_k_index[14583] = 68138;
mem_k_index[14584] = 68141;
mem_k_index[14585] = 68143;
mem_k_index[14586] = 68146;
mem_k_index[14587] = 68148;
mem_k_index[14588] = 68151;
mem_k_index[14589] = 68153;
mem_k_index[14590] = 68156;
mem_k_index[14591] = 68158;
mem_k_index[14592] = 68480;
mem_k_index[14593] = 68482;
mem_k_index[14594] = 68485;
mem_k_index[14595] = 68487;
mem_k_index[14596] = 68490;
mem_k_index[14597] = 68492;
mem_k_index[14598] = 68495;
mem_k_index[14599] = 68497;
mem_k_index[14600] = 68500;
mem_k_index[14601] = 68502;
mem_k_index[14602] = 68505;
mem_k_index[14603] = 68507;
mem_k_index[14604] = 68510;
mem_k_index[14605] = 68512;
mem_k_index[14606] = 68515;
mem_k_index[14607] = 68517;
mem_k_index[14608] = 68520;
mem_k_index[14609] = 68522;
mem_k_index[14610] = 68525;
mem_k_index[14611] = 68527;
mem_k_index[14612] = 68530;
mem_k_index[14613] = 68532;
mem_k_index[14614] = 68535;
mem_k_index[14615] = 68537;
mem_k_index[14616] = 68540;
mem_k_index[14617] = 68542;
mem_k_index[14618] = 68545;
mem_k_index[14619] = 68547;
mem_k_index[14620] = 68550;
mem_k_index[14621] = 68552;
mem_k_index[14622] = 68555;
mem_k_index[14623] = 68557;
mem_k_index[14624] = 68560;
mem_k_index[14625] = 68562;
mem_k_index[14626] = 68565;
mem_k_index[14627] = 68567;
mem_k_index[14628] = 68570;
mem_k_index[14629] = 68572;
mem_k_index[14630] = 68575;
mem_k_index[14631] = 68577;
mem_k_index[14632] = 68580;
mem_k_index[14633] = 68582;
mem_k_index[14634] = 68585;
mem_k_index[14635] = 68588;
mem_k_index[14636] = 68590;
mem_k_index[14637] = 68593;
mem_k_index[14638] = 68595;
mem_k_index[14639] = 68598;
mem_k_index[14640] = 68600;
mem_k_index[14641] = 68603;
mem_k_index[14642] = 68605;
mem_k_index[14643] = 68608;
mem_k_index[14644] = 68610;
mem_k_index[14645] = 68613;
mem_k_index[14646] = 68615;
mem_k_index[14647] = 68618;
mem_k_index[14648] = 68620;
mem_k_index[14649] = 68623;
mem_k_index[14650] = 68625;
mem_k_index[14651] = 68628;
mem_k_index[14652] = 68630;
mem_k_index[14653] = 68633;
mem_k_index[14654] = 68635;
mem_k_index[14655] = 68638;
mem_k_index[14656] = 68640;
mem_k_index[14657] = 68643;
mem_k_index[14658] = 68645;
mem_k_index[14659] = 68648;
mem_k_index[14660] = 68650;
mem_k_index[14661] = 68653;
mem_k_index[14662] = 68655;
mem_k_index[14663] = 68658;
mem_k_index[14664] = 68660;
mem_k_index[14665] = 68663;
mem_k_index[14666] = 68665;
mem_k_index[14667] = 68668;
mem_k_index[14668] = 68670;
mem_k_index[14669] = 68673;
mem_k_index[14670] = 68675;
mem_k_index[14671] = 68678;
mem_k_index[14672] = 68680;
mem_k_index[14673] = 68683;
mem_k_index[14674] = 68685;
mem_k_index[14675] = 68688;
mem_k_index[14676] = 68690;
mem_k_index[14677] = 68693;
mem_k_index[14678] = 68696;
mem_k_index[14679] = 68698;
mem_k_index[14680] = 68701;
mem_k_index[14681] = 68703;
mem_k_index[14682] = 68706;
mem_k_index[14683] = 68708;
mem_k_index[14684] = 68711;
mem_k_index[14685] = 68713;
mem_k_index[14686] = 68716;
mem_k_index[14687] = 68718;
mem_k_index[14688] = 68721;
mem_k_index[14689] = 68723;
mem_k_index[14690] = 68726;
mem_k_index[14691] = 68728;
mem_k_index[14692] = 68731;
mem_k_index[14693] = 68733;
mem_k_index[14694] = 68736;
mem_k_index[14695] = 68738;
mem_k_index[14696] = 68741;
mem_k_index[14697] = 68743;
mem_k_index[14698] = 68746;
mem_k_index[14699] = 68748;
mem_k_index[14700] = 68751;
mem_k_index[14701] = 68753;
mem_k_index[14702] = 68756;
mem_k_index[14703] = 68758;
mem_k_index[14704] = 68761;
mem_k_index[14705] = 68763;
mem_k_index[14706] = 68766;
mem_k_index[14707] = 68768;
mem_k_index[14708] = 68771;
mem_k_index[14709] = 68773;
mem_k_index[14710] = 68776;
mem_k_index[14711] = 68778;
mem_k_index[14712] = 68781;
mem_k_index[14713] = 68783;
mem_k_index[14714] = 68786;
mem_k_index[14715] = 68788;
mem_k_index[14716] = 68791;
mem_k_index[14717] = 68793;
mem_k_index[14718] = 68796;
mem_k_index[14719] = 68798;
mem_k_index[14720] = 69120;
mem_k_index[14721] = 69122;
mem_k_index[14722] = 69125;
mem_k_index[14723] = 69127;
mem_k_index[14724] = 69130;
mem_k_index[14725] = 69132;
mem_k_index[14726] = 69135;
mem_k_index[14727] = 69137;
mem_k_index[14728] = 69140;
mem_k_index[14729] = 69142;
mem_k_index[14730] = 69145;
mem_k_index[14731] = 69147;
mem_k_index[14732] = 69150;
mem_k_index[14733] = 69152;
mem_k_index[14734] = 69155;
mem_k_index[14735] = 69157;
mem_k_index[14736] = 69160;
mem_k_index[14737] = 69162;
mem_k_index[14738] = 69165;
mem_k_index[14739] = 69167;
mem_k_index[14740] = 69170;
mem_k_index[14741] = 69172;
mem_k_index[14742] = 69175;
mem_k_index[14743] = 69177;
mem_k_index[14744] = 69180;
mem_k_index[14745] = 69182;
mem_k_index[14746] = 69185;
mem_k_index[14747] = 69187;
mem_k_index[14748] = 69190;
mem_k_index[14749] = 69192;
mem_k_index[14750] = 69195;
mem_k_index[14751] = 69197;
mem_k_index[14752] = 69200;
mem_k_index[14753] = 69202;
mem_k_index[14754] = 69205;
mem_k_index[14755] = 69207;
mem_k_index[14756] = 69210;
mem_k_index[14757] = 69212;
mem_k_index[14758] = 69215;
mem_k_index[14759] = 69217;
mem_k_index[14760] = 69220;
mem_k_index[14761] = 69222;
mem_k_index[14762] = 69225;
mem_k_index[14763] = 69228;
mem_k_index[14764] = 69230;
mem_k_index[14765] = 69233;
mem_k_index[14766] = 69235;
mem_k_index[14767] = 69238;
mem_k_index[14768] = 69240;
mem_k_index[14769] = 69243;
mem_k_index[14770] = 69245;
mem_k_index[14771] = 69248;
mem_k_index[14772] = 69250;
mem_k_index[14773] = 69253;
mem_k_index[14774] = 69255;
mem_k_index[14775] = 69258;
mem_k_index[14776] = 69260;
mem_k_index[14777] = 69263;
mem_k_index[14778] = 69265;
mem_k_index[14779] = 69268;
mem_k_index[14780] = 69270;
mem_k_index[14781] = 69273;
mem_k_index[14782] = 69275;
mem_k_index[14783] = 69278;
mem_k_index[14784] = 69280;
mem_k_index[14785] = 69283;
mem_k_index[14786] = 69285;
mem_k_index[14787] = 69288;
mem_k_index[14788] = 69290;
mem_k_index[14789] = 69293;
mem_k_index[14790] = 69295;
mem_k_index[14791] = 69298;
mem_k_index[14792] = 69300;
mem_k_index[14793] = 69303;
mem_k_index[14794] = 69305;
mem_k_index[14795] = 69308;
mem_k_index[14796] = 69310;
mem_k_index[14797] = 69313;
mem_k_index[14798] = 69315;
mem_k_index[14799] = 69318;
mem_k_index[14800] = 69320;
mem_k_index[14801] = 69323;
mem_k_index[14802] = 69325;
mem_k_index[14803] = 69328;
mem_k_index[14804] = 69330;
mem_k_index[14805] = 69333;
mem_k_index[14806] = 69336;
mem_k_index[14807] = 69338;
mem_k_index[14808] = 69341;
mem_k_index[14809] = 69343;
mem_k_index[14810] = 69346;
mem_k_index[14811] = 69348;
mem_k_index[14812] = 69351;
mem_k_index[14813] = 69353;
mem_k_index[14814] = 69356;
mem_k_index[14815] = 69358;
mem_k_index[14816] = 69361;
mem_k_index[14817] = 69363;
mem_k_index[14818] = 69366;
mem_k_index[14819] = 69368;
mem_k_index[14820] = 69371;
mem_k_index[14821] = 69373;
mem_k_index[14822] = 69376;
mem_k_index[14823] = 69378;
mem_k_index[14824] = 69381;
mem_k_index[14825] = 69383;
mem_k_index[14826] = 69386;
mem_k_index[14827] = 69388;
mem_k_index[14828] = 69391;
mem_k_index[14829] = 69393;
mem_k_index[14830] = 69396;
mem_k_index[14831] = 69398;
mem_k_index[14832] = 69401;
mem_k_index[14833] = 69403;
mem_k_index[14834] = 69406;
mem_k_index[14835] = 69408;
mem_k_index[14836] = 69411;
mem_k_index[14837] = 69413;
mem_k_index[14838] = 69416;
mem_k_index[14839] = 69418;
mem_k_index[14840] = 69421;
mem_k_index[14841] = 69423;
mem_k_index[14842] = 69426;
mem_k_index[14843] = 69428;
mem_k_index[14844] = 69431;
mem_k_index[14845] = 69433;
mem_k_index[14846] = 69436;
mem_k_index[14847] = 69438;
mem_k_index[14848] = 69760;
mem_k_index[14849] = 69762;
mem_k_index[14850] = 69765;
mem_k_index[14851] = 69767;
mem_k_index[14852] = 69770;
mem_k_index[14853] = 69772;
mem_k_index[14854] = 69775;
mem_k_index[14855] = 69777;
mem_k_index[14856] = 69780;
mem_k_index[14857] = 69782;
mem_k_index[14858] = 69785;
mem_k_index[14859] = 69787;
mem_k_index[14860] = 69790;
mem_k_index[14861] = 69792;
mem_k_index[14862] = 69795;
mem_k_index[14863] = 69797;
mem_k_index[14864] = 69800;
mem_k_index[14865] = 69802;
mem_k_index[14866] = 69805;
mem_k_index[14867] = 69807;
mem_k_index[14868] = 69810;
mem_k_index[14869] = 69812;
mem_k_index[14870] = 69815;
mem_k_index[14871] = 69817;
mem_k_index[14872] = 69820;
mem_k_index[14873] = 69822;
mem_k_index[14874] = 69825;
mem_k_index[14875] = 69827;
mem_k_index[14876] = 69830;
mem_k_index[14877] = 69832;
mem_k_index[14878] = 69835;
mem_k_index[14879] = 69837;
mem_k_index[14880] = 69840;
mem_k_index[14881] = 69842;
mem_k_index[14882] = 69845;
mem_k_index[14883] = 69847;
mem_k_index[14884] = 69850;
mem_k_index[14885] = 69852;
mem_k_index[14886] = 69855;
mem_k_index[14887] = 69857;
mem_k_index[14888] = 69860;
mem_k_index[14889] = 69862;
mem_k_index[14890] = 69865;
mem_k_index[14891] = 69868;
mem_k_index[14892] = 69870;
mem_k_index[14893] = 69873;
mem_k_index[14894] = 69875;
mem_k_index[14895] = 69878;
mem_k_index[14896] = 69880;
mem_k_index[14897] = 69883;
mem_k_index[14898] = 69885;
mem_k_index[14899] = 69888;
mem_k_index[14900] = 69890;
mem_k_index[14901] = 69893;
mem_k_index[14902] = 69895;
mem_k_index[14903] = 69898;
mem_k_index[14904] = 69900;
mem_k_index[14905] = 69903;
mem_k_index[14906] = 69905;
mem_k_index[14907] = 69908;
mem_k_index[14908] = 69910;
mem_k_index[14909] = 69913;
mem_k_index[14910] = 69915;
mem_k_index[14911] = 69918;
mem_k_index[14912] = 69920;
mem_k_index[14913] = 69923;
mem_k_index[14914] = 69925;
mem_k_index[14915] = 69928;
mem_k_index[14916] = 69930;
mem_k_index[14917] = 69933;
mem_k_index[14918] = 69935;
mem_k_index[14919] = 69938;
mem_k_index[14920] = 69940;
mem_k_index[14921] = 69943;
mem_k_index[14922] = 69945;
mem_k_index[14923] = 69948;
mem_k_index[14924] = 69950;
mem_k_index[14925] = 69953;
mem_k_index[14926] = 69955;
mem_k_index[14927] = 69958;
mem_k_index[14928] = 69960;
mem_k_index[14929] = 69963;
mem_k_index[14930] = 69965;
mem_k_index[14931] = 69968;
mem_k_index[14932] = 69970;
mem_k_index[14933] = 69973;
mem_k_index[14934] = 69976;
mem_k_index[14935] = 69978;
mem_k_index[14936] = 69981;
mem_k_index[14937] = 69983;
mem_k_index[14938] = 69986;
mem_k_index[14939] = 69988;
mem_k_index[14940] = 69991;
mem_k_index[14941] = 69993;
mem_k_index[14942] = 69996;
mem_k_index[14943] = 69998;
mem_k_index[14944] = 70001;
mem_k_index[14945] = 70003;
mem_k_index[14946] = 70006;
mem_k_index[14947] = 70008;
mem_k_index[14948] = 70011;
mem_k_index[14949] = 70013;
mem_k_index[14950] = 70016;
mem_k_index[14951] = 70018;
mem_k_index[14952] = 70021;
mem_k_index[14953] = 70023;
mem_k_index[14954] = 70026;
mem_k_index[14955] = 70028;
mem_k_index[14956] = 70031;
mem_k_index[14957] = 70033;
mem_k_index[14958] = 70036;
mem_k_index[14959] = 70038;
mem_k_index[14960] = 70041;
mem_k_index[14961] = 70043;
mem_k_index[14962] = 70046;
mem_k_index[14963] = 70048;
mem_k_index[14964] = 70051;
mem_k_index[14965] = 70053;
mem_k_index[14966] = 70056;
mem_k_index[14967] = 70058;
mem_k_index[14968] = 70061;
mem_k_index[14969] = 70063;
mem_k_index[14970] = 70066;
mem_k_index[14971] = 70068;
mem_k_index[14972] = 70071;
mem_k_index[14973] = 70073;
mem_k_index[14974] = 70076;
mem_k_index[14975] = 70078;
mem_k_index[14976] = 70400;
mem_k_index[14977] = 70402;
mem_k_index[14978] = 70405;
mem_k_index[14979] = 70407;
mem_k_index[14980] = 70410;
mem_k_index[14981] = 70412;
mem_k_index[14982] = 70415;
mem_k_index[14983] = 70417;
mem_k_index[14984] = 70420;
mem_k_index[14985] = 70422;
mem_k_index[14986] = 70425;
mem_k_index[14987] = 70427;
mem_k_index[14988] = 70430;
mem_k_index[14989] = 70432;
mem_k_index[14990] = 70435;
mem_k_index[14991] = 70437;
mem_k_index[14992] = 70440;
mem_k_index[14993] = 70442;
mem_k_index[14994] = 70445;
mem_k_index[14995] = 70447;
mem_k_index[14996] = 70450;
mem_k_index[14997] = 70452;
mem_k_index[14998] = 70455;
mem_k_index[14999] = 70457;
mem_k_index[15000] = 70460;
mem_k_index[15001] = 70462;
mem_k_index[15002] = 70465;
mem_k_index[15003] = 70467;
mem_k_index[15004] = 70470;
mem_k_index[15005] = 70472;
mem_k_index[15006] = 70475;
mem_k_index[15007] = 70477;
mem_k_index[15008] = 70480;
mem_k_index[15009] = 70482;
mem_k_index[15010] = 70485;
mem_k_index[15011] = 70487;
mem_k_index[15012] = 70490;
mem_k_index[15013] = 70492;
mem_k_index[15014] = 70495;
mem_k_index[15015] = 70497;
mem_k_index[15016] = 70500;
mem_k_index[15017] = 70502;
mem_k_index[15018] = 70505;
mem_k_index[15019] = 70508;
mem_k_index[15020] = 70510;
mem_k_index[15021] = 70513;
mem_k_index[15022] = 70515;
mem_k_index[15023] = 70518;
mem_k_index[15024] = 70520;
mem_k_index[15025] = 70523;
mem_k_index[15026] = 70525;
mem_k_index[15027] = 70528;
mem_k_index[15028] = 70530;
mem_k_index[15029] = 70533;
mem_k_index[15030] = 70535;
mem_k_index[15031] = 70538;
mem_k_index[15032] = 70540;
mem_k_index[15033] = 70543;
mem_k_index[15034] = 70545;
mem_k_index[15035] = 70548;
mem_k_index[15036] = 70550;
mem_k_index[15037] = 70553;
mem_k_index[15038] = 70555;
mem_k_index[15039] = 70558;
mem_k_index[15040] = 70560;
mem_k_index[15041] = 70563;
mem_k_index[15042] = 70565;
mem_k_index[15043] = 70568;
mem_k_index[15044] = 70570;
mem_k_index[15045] = 70573;
mem_k_index[15046] = 70575;
mem_k_index[15047] = 70578;
mem_k_index[15048] = 70580;
mem_k_index[15049] = 70583;
mem_k_index[15050] = 70585;
mem_k_index[15051] = 70588;
mem_k_index[15052] = 70590;
mem_k_index[15053] = 70593;
mem_k_index[15054] = 70595;
mem_k_index[15055] = 70598;
mem_k_index[15056] = 70600;
mem_k_index[15057] = 70603;
mem_k_index[15058] = 70605;
mem_k_index[15059] = 70608;
mem_k_index[15060] = 70610;
mem_k_index[15061] = 70613;
mem_k_index[15062] = 70616;
mem_k_index[15063] = 70618;
mem_k_index[15064] = 70621;
mem_k_index[15065] = 70623;
mem_k_index[15066] = 70626;
mem_k_index[15067] = 70628;
mem_k_index[15068] = 70631;
mem_k_index[15069] = 70633;
mem_k_index[15070] = 70636;
mem_k_index[15071] = 70638;
mem_k_index[15072] = 70641;
mem_k_index[15073] = 70643;
mem_k_index[15074] = 70646;
mem_k_index[15075] = 70648;
mem_k_index[15076] = 70651;
mem_k_index[15077] = 70653;
mem_k_index[15078] = 70656;
mem_k_index[15079] = 70658;
mem_k_index[15080] = 70661;
mem_k_index[15081] = 70663;
mem_k_index[15082] = 70666;
mem_k_index[15083] = 70668;
mem_k_index[15084] = 70671;
mem_k_index[15085] = 70673;
mem_k_index[15086] = 70676;
mem_k_index[15087] = 70678;
mem_k_index[15088] = 70681;
mem_k_index[15089] = 70683;
mem_k_index[15090] = 70686;
mem_k_index[15091] = 70688;
mem_k_index[15092] = 70691;
mem_k_index[15093] = 70693;
mem_k_index[15094] = 70696;
mem_k_index[15095] = 70698;
mem_k_index[15096] = 70701;
mem_k_index[15097] = 70703;
mem_k_index[15098] = 70706;
mem_k_index[15099] = 70708;
mem_k_index[15100] = 70711;
mem_k_index[15101] = 70713;
mem_k_index[15102] = 70716;
mem_k_index[15103] = 70718;
mem_k_index[15104] = 71040;
mem_k_index[15105] = 71042;
mem_k_index[15106] = 71045;
mem_k_index[15107] = 71047;
mem_k_index[15108] = 71050;
mem_k_index[15109] = 71052;
mem_k_index[15110] = 71055;
mem_k_index[15111] = 71057;
mem_k_index[15112] = 71060;
mem_k_index[15113] = 71062;
mem_k_index[15114] = 71065;
mem_k_index[15115] = 71067;
mem_k_index[15116] = 71070;
mem_k_index[15117] = 71072;
mem_k_index[15118] = 71075;
mem_k_index[15119] = 71077;
mem_k_index[15120] = 71080;
mem_k_index[15121] = 71082;
mem_k_index[15122] = 71085;
mem_k_index[15123] = 71087;
mem_k_index[15124] = 71090;
mem_k_index[15125] = 71092;
mem_k_index[15126] = 71095;
mem_k_index[15127] = 71097;
mem_k_index[15128] = 71100;
mem_k_index[15129] = 71102;
mem_k_index[15130] = 71105;
mem_k_index[15131] = 71107;
mem_k_index[15132] = 71110;
mem_k_index[15133] = 71112;
mem_k_index[15134] = 71115;
mem_k_index[15135] = 71117;
mem_k_index[15136] = 71120;
mem_k_index[15137] = 71122;
mem_k_index[15138] = 71125;
mem_k_index[15139] = 71127;
mem_k_index[15140] = 71130;
mem_k_index[15141] = 71132;
mem_k_index[15142] = 71135;
mem_k_index[15143] = 71137;
mem_k_index[15144] = 71140;
mem_k_index[15145] = 71142;
mem_k_index[15146] = 71145;
mem_k_index[15147] = 71148;
mem_k_index[15148] = 71150;
mem_k_index[15149] = 71153;
mem_k_index[15150] = 71155;
mem_k_index[15151] = 71158;
mem_k_index[15152] = 71160;
mem_k_index[15153] = 71163;
mem_k_index[15154] = 71165;
mem_k_index[15155] = 71168;
mem_k_index[15156] = 71170;
mem_k_index[15157] = 71173;
mem_k_index[15158] = 71175;
mem_k_index[15159] = 71178;
mem_k_index[15160] = 71180;
mem_k_index[15161] = 71183;
mem_k_index[15162] = 71185;
mem_k_index[15163] = 71188;
mem_k_index[15164] = 71190;
mem_k_index[15165] = 71193;
mem_k_index[15166] = 71195;
mem_k_index[15167] = 71198;
mem_k_index[15168] = 71200;
mem_k_index[15169] = 71203;
mem_k_index[15170] = 71205;
mem_k_index[15171] = 71208;
mem_k_index[15172] = 71210;
mem_k_index[15173] = 71213;
mem_k_index[15174] = 71215;
mem_k_index[15175] = 71218;
mem_k_index[15176] = 71220;
mem_k_index[15177] = 71223;
mem_k_index[15178] = 71225;
mem_k_index[15179] = 71228;
mem_k_index[15180] = 71230;
mem_k_index[15181] = 71233;
mem_k_index[15182] = 71235;
mem_k_index[15183] = 71238;
mem_k_index[15184] = 71240;
mem_k_index[15185] = 71243;
mem_k_index[15186] = 71245;
mem_k_index[15187] = 71248;
mem_k_index[15188] = 71250;
mem_k_index[15189] = 71253;
mem_k_index[15190] = 71256;
mem_k_index[15191] = 71258;
mem_k_index[15192] = 71261;
mem_k_index[15193] = 71263;
mem_k_index[15194] = 71266;
mem_k_index[15195] = 71268;
mem_k_index[15196] = 71271;
mem_k_index[15197] = 71273;
mem_k_index[15198] = 71276;
mem_k_index[15199] = 71278;
mem_k_index[15200] = 71281;
mem_k_index[15201] = 71283;
mem_k_index[15202] = 71286;
mem_k_index[15203] = 71288;
mem_k_index[15204] = 71291;
mem_k_index[15205] = 71293;
mem_k_index[15206] = 71296;
mem_k_index[15207] = 71298;
mem_k_index[15208] = 71301;
mem_k_index[15209] = 71303;
mem_k_index[15210] = 71306;
mem_k_index[15211] = 71308;
mem_k_index[15212] = 71311;
mem_k_index[15213] = 71313;
mem_k_index[15214] = 71316;
mem_k_index[15215] = 71318;
mem_k_index[15216] = 71321;
mem_k_index[15217] = 71323;
mem_k_index[15218] = 71326;
mem_k_index[15219] = 71328;
mem_k_index[15220] = 71331;
mem_k_index[15221] = 71333;
mem_k_index[15222] = 71336;
mem_k_index[15223] = 71338;
mem_k_index[15224] = 71341;
mem_k_index[15225] = 71343;
mem_k_index[15226] = 71346;
mem_k_index[15227] = 71348;
mem_k_index[15228] = 71351;
mem_k_index[15229] = 71353;
mem_k_index[15230] = 71356;
mem_k_index[15231] = 71358;
mem_k_index[15232] = 71360;
mem_k_index[15233] = 71362;
mem_k_index[15234] = 71365;
mem_k_index[15235] = 71367;
mem_k_index[15236] = 71370;
mem_k_index[15237] = 71372;
mem_k_index[15238] = 71375;
mem_k_index[15239] = 71377;
mem_k_index[15240] = 71380;
mem_k_index[15241] = 71382;
mem_k_index[15242] = 71385;
mem_k_index[15243] = 71387;
mem_k_index[15244] = 71390;
mem_k_index[15245] = 71392;
mem_k_index[15246] = 71395;
mem_k_index[15247] = 71397;
mem_k_index[15248] = 71400;
mem_k_index[15249] = 71402;
mem_k_index[15250] = 71405;
mem_k_index[15251] = 71407;
mem_k_index[15252] = 71410;
mem_k_index[15253] = 71412;
mem_k_index[15254] = 71415;
mem_k_index[15255] = 71417;
mem_k_index[15256] = 71420;
mem_k_index[15257] = 71422;
mem_k_index[15258] = 71425;
mem_k_index[15259] = 71427;
mem_k_index[15260] = 71430;
mem_k_index[15261] = 71432;
mem_k_index[15262] = 71435;
mem_k_index[15263] = 71437;
mem_k_index[15264] = 71440;
mem_k_index[15265] = 71442;
mem_k_index[15266] = 71445;
mem_k_index[15267] = 71447;
mem_k_index[15268] = 71450;
mem_k_index[15269] = 71452;
mem_k_index[15270] = 71455;
mem_k_index[15271] = 71457;
mem_k_index[15272] = 71460;
mem_k_index[15273] = 71462;
mem_k_index[15274] = 71465;
mem_k_index[15275] = 71468;
mem_k_index[15276] = 71470;
mem_k_index[15277] = 71473;
mem_k_index[15278] = 71475;
mem_k_index[15279] = 71478;
mem_k_index[15280] = 71480;
mem_k_index[15281] = 71483;
mem_k_index[15282] = 71485;
mem_k_index[15283] = 71488;
mem_k_index[15284] = 71490;
mem_k_index[15285] = 71493;
mem_k_index[15286] = 71495;
mem_k_index[15287] = 71498;
mem_k_index[15288] = 71500;
mem_k_index[15289] = 71503;
mem_k_index[15290] = 71505;
mem_k_index[15291] = 71508;
mem_k_index[15292] = 71510;
mem_k_index[15293] = 71513;
mem_k_index[15294] = 71515;
mem_k_index[15295] = 71518;
mem_k_index[15296] = 71520;
mem_k_index[15297] = 71523;
mem_k_index[15298] = 71525;
mem_k_index[15299] = 71528;
mem_k_index[15300] = 71530;
mem_k_index[15301] = 71533;
mem_k_index[15302] = 71535;
mem_k_index[15303] = 71538;
mem_k_index[15304] = 71540;
mem_k_index[15305] = 71543;
mem_k_index[15306] = 71545;
mem_k_index[15307] = 71548;
mem_k_index[15308] = 71550;
mem_k_index[15309] = 71553;
mem_k_index[15310] = 71555;
mem_k_index[15311] = 71558;
mem_k_index[15312] = 71560;
mem_k_index[15313] = 71563;
mem_k_index[15314] = 71565;
mem_k_index[15315] = 71568;
mem_k_index[15316] = 71570;
mem_k_index[15317] = 71573;
mem_k_index[15318] = 71576;
mem_k_index[15319] = 71578;
mem_k_index[15320] = 71581;
mem_k_index[15321] = 71583;
mem_k_index[15322] = 71586;
mem_k_index[15323] = 71588;
mem_k_index[15324] = 71591;
mem_k_index[15325] = 71593;
mem_k_index[15326] = 71596;
mem_k_index[15327] = 71598;
mem_k_index[15328] = 71601;
mem_k_index[15329] = 71603;
mem_k_index[15330] = 71606;
mem_k_index[15331] = 71608;
mem_k_index[15332] = 71611;
mem_k_index[15333] = 71613;
mem_k_index[15334] = 71616;
mem_k_index[15335] = 71618;
mem_k_index[15336] = 71621;
mem_k_index[15337] = 71623;
mem_k_index[15338] = 71626;
mem_k_index[15339] = 71628;
mem_k_index[15340] = 71631;
mem_k_index[15341] = 71633;
mem_k_index[15342] = 71636;
mem_k_index[15343] = 71638;
mem_k_index[15344] = 71641;
mem_k_index[15345] = 71643;
mem_k_index[15346] = 71646;
mem_k_index[15347] = 71648;
mem_k_index[15348] = 71651;
mem_k_index[15349] = 71653;
mem_k_index[15350] = 71656;
mem_k_index[15351] = 71658;
mem_k_index[15352] = 71661;
mem_k_index[15353] = 71663;
mem_k_index[15354] = 71666;
mem_k_index[15355] = 71668;
mem_k_index[15356] = 71671;
mem_k_index[15357] = 71673;
mem_k_index[15358] = 71676;
mem_k_index[15359] = 71678;
mem_k_index[15360] = 72000;
mem_k_index[15361] = 72002;
mem_k_index[15362] = 72005;
mem_k_index[15363] = 72007;
mem_k_index[15364] = 72010;
mem_k_index[15365] = 72012;
mem_k_index[15366] = 72015;
mem_k_index[15367] = 72017;
mem_k_index[15368] = 72020;
mem_k_index[15369] = 72022;
mem_k_index[15370] = 72025;
mem_k_index[15371] = 72027;
mem_k_index[15372] = 72030;
mem_k_index[15373] = 72032;
mem_k_index[15374] = 72035;
mem_k_index[15375] = 72037;
mem_k_index[15376] = 72040;
mem_k_index[15377] = 72042;
mem_k_index[15378] = 72045;
mem_k_index[15379] = 72047;
mem_k_index[15380] = 72050;
mem_k_index[15381] = 72052;
mem_k_index[15382] = 72055;
mem_k_index[15383] = 72057;
mem_k_index[15384] = 72060;
mem_k_index[15385] = 72062;
mem_k_index[15386] = 72065;
mem_k_index[15387] = 72067;
mem_k_index[15388] = 72070;
mem_k_index[15389] = 72072;
mem_k_index[15390] = 72075;
mem_k_index[15391] = 72077;
mem_k_index[15392] = 72080;
mem_k_index[15393] = 72082;
mem_k_index[15394] = 72085;
mem_k_index[15395] = 72087;
mem_k_index[15396] = 72090;
mem_k_index[15397] = 72092;
mem_k_index[15398] = 72095;
mem_k_index[15399] = 72097;
mem_k_index[15400] = 72100;
mem_k_index[15401] = 72102;
mem_k_index[15402] = 72105;
mem_k_index[15403] = 72108;
mem_k_index[15404] = 72110;
mem_k_index[15405] = 72113;
mem_k_index[15406] = 72115;
mem_k_index[15407] = 72118;
mem_k_index[15408] = 72120;
mem_k_index[15409] = 72123;
mem_k_index[15410] = 72125;
mem_k_index[15411] = 72128;
mem_k_index[15412] = 72130;
mem_k_index[15413] = 72133;
mem_k_index[15414] = 72135;
mem_k_index[15415] = 72138;
mem_k_index[15416] = 72140;
mem_k_index[15417] = 72143;
mem_k_index[15418] = 72145;
mem_k_index[15419] = 72148;
mem_k_index[15420] = 72150;
mem_k_index[15421] = 72153;
mem_k_index[15422] = 72155;
mem_k_index[15423] = 72158;
mem_k_index[15424] = 72160;
mem_k_index[15425] = 72163;
mem_k_index[15426] = 72165;
mem_k_index[15427] = 72168;
mem_k_index[15428] = 72170;
mem_k_index[15429] = 72173;
mem_k_index[15430] = 72175;
mem_k_index[15431] = 72178;
mem_k_index[15432] = 72180;
mem_k_index[15433] = 72183;
mem_k_index[15434] = 72185;
mem_k_index[15435] = 72188;
mem_k_index[15436] = 72190;
mem_k_index[15437] = 72193;
mem_k_index[15438] = 72195;
mem_k_index[15439] = 72198;
mem_k_index[15440] = 72200;
mem_k_index[15441] = 72203;
mem_k_index[15442] = 72205;
mem_k_index[15443] = 72208;
mem_k_index[15444] = 72210;
mem_k_index[15445] = 72213;
mem_k_index[15446] = 72216;
mem_k_index[15447] = 72218;
mem_k_index[15448] = 72221;
mem_k_index[15449] = 72223;
mem_k_index[15450] = 72226;
mem_k_index[15451] = 72228;
mem_k_index[15452] = 72231;
mem_k_index[15453] = 72233;
mem_k_index[15454] = 72236;
mem_k_index[15455] = 72238;
mem_k_index[15456] = 72241;
mem_k_index[15457] = 72243;
mem_k_index[15458] = 72246;
mem_k_index[15459] = 72248;
mem_k_index[15460] = 72251;
mem_k_index[15461] = 72253;
mem_k_index[15462] = 72256;
mem_k_index[15463] = 72258;
mem_k_index[15464] = 72261;
mem_k_index[15465] = 72263;
mem_k_index[15466] = 72266;
mem_k_index[15467] = 72268;
mem_k_index[15468] = 72271;
mem_k_index[15469] = 72273;
mem_k_index[15470] = 72276;
mem_k_index[15471] = 72278;
mem_k_index[15472] = 72281;
mem_k_index[15473] = 72283;
mem_k_index[15474] = 72286;
mem_k_index[15475] = 72288;
mem_k_index[15476] = 72291;
mem_k_index[15477] = 72293;
mem_k_index[15478] = 72296;
mem_k_index[15479] = 72298;
mem_k_index[15480] = 72301;
mem_k_index[15481] = 72303;
mem_k_index[15482] = 72306;
mem_k_index[15483] = 72308;
mem_k_index[15484] = 72311;
mem_k_index[15485] = 72313;
mem_k_index[15486] = 72316;
mem_k_index[15487] = 72318;
mem_k_index[15488] = 72640;
mem_k_index[15489] = 72642;
mem_k_index[15490] = 72645;
mem_k_index[15491] = 72647;
mem_k_index[15492] = 72650;
mem_k_index[15493] = 72652;
mem_k_index[15494] = 72655;
mem_k_index[15495] = 72657;
mem_k_index[15496] = 72660;
mem_k_index[15497] = 72662;
mem_k_index[15498] = 72665;
mem_k_index[15499] = 72667;
mem_k_index[15500] = 72670;
mem_k_index[15501] = 72672;
mem_k_index[15502] = 72675;
mem_k_index[15503] = 72677;
mem_k_index[15504] = 72680;
mem_k_index[15505] = 72682;
mem_k_index[15506] = 72685;
mem_k_index[15507] = 72687;
mem_k_index[15508] = 72690;
mem_k_index[15509] = 72692;
mem_k_index[15510] = 72695;
mem_k_index[15511] = 72697;
mem_k_index[15512] = 72700;
mem_k_index[15513] = 72702;
mem_k_index[15514] = 72705;
mem_k_index[15515] = 72707;
mem_k_index[15516] = 72710;
mem_k_index[15517] = 72712;
mem_k_index[15518] = 72715;
mem_k_index[15519] = 72717;
mem_k_index[15520] = 72720;
mem_k_index[15521] = 72722;
mem_k_index[15522] = 72725;
mem_k_index[15523] = 72727;
mem_k_index[15524] = 72730;
mem_k_index[15525] = 72732;
mem_k_index[15526] = 72735;
mem_k_index[15527] = 72737;
mem_k_index[15528] = 72740;
mem_k_index[15529] = 72742;
mem_k_index[15530] = 72745;
mem_k_index[15531] = 72748;
mem_k_index[15532] = 72750;
mem_k_index[15533] = 72753;
mem_k_index[15534] = 72755;
mem_k_index[15535] = 72758;
mem_k_index[15536] = 72760;
mem_k_index[15537] = 72763;
mem_k_index[15538] = 72765;
mem_k_index[15539] = 72768;
mem_k_index[15540] = 72770;
mem_k_index[15541] = 72773;
mem_k_index[15542] = 72775;
mem_k_index[15543] = 72778;
mem_k_index[15544] = 72780;
mem_k_index[15545] = 72783;
mem_k_index[15546] = 72785;
mem_k_index[15547] = 72788;
mem_k_index[15548] = 72790;
mem_k_index[15549] = 72793;
mem_k_index[15550] = 72795;
mem_k_index[15551] = 72798;
mem_k_index[15552] = 72800;
mem_k_index[15553] = 72803;
mem_k_index[15554] = 72805;
mem_k_index[15555] = 72808;
mem_k_index[15556] = 72810;
mem_k_index[15557] = 72813;
mem_k_index[15558] = 72815;
mem_k_index[15559] = 72818;
mem_k_index[15560] = 72820;
mem_k_index[15561] = 72823;
mem_k_index[15562] = 72825;
mem_k_index[15563] = 72828;
mem_k_index[15564] = 72830;
mem_k_index[15565] = 72833;
mem_k_index[15566] = 72835;
mem_k_index[15567] = 72838;
mem_k_index[15568] = 72840;
mem_k_index[15569] = 72843;
mem_k_index[15570] = 72845;
mem_k_index[15571] = 72848;
mem_k_index[15572] = 72850;
mem_k_index[15573] = 72853;
mem_k_index[15574] = 72856;
mem_k_index[15575] = 72858;
mem_k_index[15576] = 72861;
mem_k_index[15577] = 72863;
mem_k_index[15578] = 72866;
mem_k_index[15579] = 72868;
mem_k_index[15580] = 72871;
mem_k_index[15581] = 72873;
mem_k_index[15582] = 72876;
mem_k_index[15583] = 72878;
mem_k_index[15584] = 72881;
mem_k_index[15585] = 72883;
mem_k_index[15586] = 72886;
mem_k_index[15587] = 72888;
mem_k_index[15588] = 72891;
mem_k_index[15589] = 72893;
mem_k_index[15590] = 72896;
mem_k_index[15591] = 72898;
mem_k_index[15592] = 72901;
mem_k_index[15593] = 72903;
mem_k_index[15594] = 72906;
mem_k_index[15595] = 72908;
mem_k_index[15596] = 72911;
mem_k_index[15597] = 72913;
mem_k_index[15598] = 72916;
mem_k_index[15599] = 72918;
mem_k_index[15600] = 72921;
mem_k_index[15601] = 72923;
mem_k_index[15602] = 72926;
mem_k_index[15603] = 72928;
mem_k_index[15604] = 72931;
mem_k_index[15605] = 72933;
mem_k_index[15606] = 72936;
mem_k_index[15607] = 72938;
mem_k_index[15608] = 72941;
mem_k_index[15609] = 72943;
mem_k_index[15610] = 72946;
mem_k_index[15611] = 72948;
mem_k_index[15612] = 72951;
mem_k_index[15613] = 72953;
mem_k_index[15614] = 72956;
mem_k_index[15615] = 72958;
mem_k_index[15616] = 73280;
mem_k_index[15617] = 73282;
mem_k_index[15618] = 73285;
mem_k_index[15619] = 73287;
mem_k_index[15620] = 73290;
mem_k_index[15621] = 73292;
mem_k_index[15622] = 73295;
mem_k_index[15623] = 73297;
mem_k_index[15624] = 73300;
mem_k_index[15625] = 73302;
mem_k_index[15626] = 73305;
mem_k_index[15627] = 73307;
mem_k_index[15628] = 73310;
mem_k_index[15629] = 73312;
mem_k_index[15630] = 73315;
mem_k_index[15631] = 73317;
mem_k_index[15632] = 73320;
mem_k_index[15633] = 73322;
mem_k_index[15634] = 73325;
mem_k_index[15635] = 73327;
mem_k_index[15636] = 73330;
mem_k_index[15637] = 73332;
mem_k_index[15638] = 73335;
mem_k_index[15639] = 73337;
mem_k_index[15640] = 73340;
mem_k_index[15641] = 73342;
mem_k_index[15642] = 73345;
mem_k_index[15643] = 73347;
mem_k_index[15644] = 73350;
mem_k_index[15645] = 73352;
mem_k_index[15646] = 73355;
mem_k_index[15647] = 73357;
mem_k_index[15648] = 73360;
mem_k_index[15649] = 73362;
mem_k_index[15650] = 73365;
mem_k_index[15651] = 73367;
mem_k_index[15652] = 73370;
mem_k_index[15653] = 73372;
mem_k_index[15654] = 73375;
mem_k_index[15655] = 73377;
mem_k_index[15656] = 73380;
mem_k_index[15657] = 73382;
mem_k_index[15658] = 73385;
mem_k_index[15659] = 73388;
mem_k_index[15660] = 73390;
mem_k_index[15661] = 73393;
mem_k_index[15662] = 73395;
mem_k_index[15663] = 73398;
mem_k_index[15664] = 73400;
mem_k_index[15665] = 73403;
mem_k_index[15666] = 73405;
mem_k_index[15667] = 73408;
mem_k_index[15668] = 73410;
mem_k_index[15669] = 73413;
mem_k_index[15670] = 73415;
mem_k_index[15671] = 73418;
mem_k_index[15672] = 73420;
mem_k_index[15673] = 73423;
mem_k_index[15674] = 73425;
mem_k_index[15675] = 73428;
mem_k_index[15676] = 73430;
mem_k_index[15677] = 73433;
mem_k_index[15678] = 73435;
mem_k_index[15679] = 73438;
mem_k_index[15680] = 73440;
mem_k_index[15681] = 73443;
mem_k_index[15682] = 73445;
mem_k_index[15683] = 73448;
mem_k_index[15684] = 73450;
mem_k_index[15685] = 73453;
mem_k_index[15686] = 73455;
mem_k_index[15687] = 73458;
mem_k_index[15688] = 73460;
mem_k_index[15689] = 73463;
mem_k_index[15690] = 73465;
mem_k_index[15691] = 73468;
mem_k_index[15692] = 73470;
mem_k_index[15693] = 73473;
mem_k_index[15694] = 73475;
mem_k_index[15695] = 73478;
mem_k_index[15696] = 73480;
mem_k_index[15697] = 73483;
mem_k_index[15698] = 73485;
mem_k_index[15699] = 73488;
mem_k_index[15700] = 73490;
mem_k_index[15701] = 73493;
mem_k_index[15702] = 73496;
mem_k_index[15703] = 73498;
mem_k_index[15704] = 73501;
mem_k_index[15705] = 73503;
mem_k_index[15706] = 73506;
mem_k_index[15707] = 73508;
mem_k_index[15708] = 73511;
mem_k_index[15709] = 73513;
mem_k_index[15710] = 73516;
mem_k_index[15711] = 73518;
mem_k_index[15712] = 73521;
mem_k_index[15713] = 73523;
mem_k_index[15714] = 73526;
mem_k_index[15715] = 73528;
mem_k_index[15716] = 73531;
mem_k_index[15717] = 73533;
mem_k_index[15718] = 73536;
mem_k_index[15719] = 73538;
mem_k_index[15720] = 73541;
mem_k_index[15721] = 73543;
mem_k_index[15722] = 73546;
mem_k_index[15723] = 73548;
mem_k_index[15724] = 73551;
mem_k_index[15725] = 73553;
mem_k_index[15726] = 73556;
mem_k_index[15727] = 73558;
mem_k_index[15728] = 73561;
mem_k_index[15729] = 73563;
mem_k_index[15730] = 73566;
mem_k_index[15731] = 73568;
mem_k_index[15732] = 73571;
mem_k_index[15733] = 73573;
mem_k_index[15734] = 73576;
mem_k_index[15735] = 73578;
mem_k_index[15736] = 73581;
mem_k_index[15737] = 73583;
mem_k_index[15738] = 73586;
mem_k_index[15739] = 73588;
mem_k_index[15740] = 73591;
mem_k_index[15741] = 73593;
mem_k_index[15742] = 73596;
mem_k_index[15743] = 73598;
mem_k_index[15744] = 73920;
mem_k_index[15745] = 73922;
mem_k_index[15746] = 73925;
mem_k_index[15747] = 73927;
mem_k_index[15748] = 73930;
mem_k_index[15749] = 73932;
mem_k_index[15750] = 73935;
mem_k_index[15751] = 73937;
mem_k_index[15752] = 73940;
mem_k_index[15753] = 73942;
mem_k_index[15754] = 73945;
mem_k_index[15755] = 73947;
mem_k_index[15756] = 73950;
mem_k_index[15757] = 73952;
mem_k_index[15758] = 73955;
mem_k_index[15759] = 73957;
mem_k_index[15760] = 73960;
mem_k_index[15761] = 73962;
mem_k_index[15762] = 73965;
mem_k_index[15763] = 73967;
mem_k_index[15764] = 73970;
mem_k_index[15765] = 73972;
mem_k_index[15766] = 73975;
mem_k_index[15767] = 73977;
mem_k_index[15768] = 73980;
mem_k_index[15769] = 73982;
mem_k_index[15770] = 73985;
mem_k_index[15771] = 73987;
mem_k_index[15772] = 73990;
mem_k_index[15773] = 73992;
mem_k_index[15774] = 73995;
mem_k_index[15775] = 73997;
mem_k_index[15776] = 74000;
mem_k_index[15777] = 74002;
mem_k_index[15778] = 74005;
mem_k_index[15779] = 74007;
mem_k_index[15780] = 74010;
mem_k_index[15781] = 74012;
mem_k_index[15782] = 74015;
mem_k_index[15783] = 74017;
mem_k_index[15784] = 74020;
mem_k_index[15785] = 74022;
mem_k_index[15786] = 74025;
mem_k_index[15787] = 74028;
mem_k_index[15788] = 74030;
mem_k_index[15789] = 74033;
mem_k_index[15790] = 74035;
mem_k_index[15791] = 74038;
mem_k_index[15792] = 74040;
mem_k_index[15793] = 74043;
mem_k_index[15794] = 74045;
mem_k_index[15795] = 74048;
mem_k_index[15796] = 74050;
mem_k_index[15797] = 74053;
mem_k_index[15798] = 74055;
mem_k_index[15799] = 74058;
mem_k_index[15800] = 74060;
mem_k_index[15801] = 74063;
mem_k_index[15802] = 74065;
mem_k_index[15803] = 74068;
mem_k_index[15804] = 74070;
mem_k_index[15805] = 74073;
mem_k_index[15806] = 74075;
mem_k_index[15807] = 74078;
mem_k_index[15808] = 74080;
mem_k_index[15809] = 74083;
mem_k_index[15810] = 74085;
mem_k_index[15811] = 74088;
mem_k_index[15812] = 74090;
mem_k_index[15813] = 74093;
mem_k_index[15814] = 74095;
mem_k_index[15815] = 74098;
mem_k_index[15816] = 74100;
mem_k_index[15817] = 74103;
mem_k_index[15818] = 74105;
mem_k_index[15819] = 74108;
mem_k_index[15820] = 74110;
mem_k_index[15821] = 74113;
mem_k_index[15822] = 74115;
mem_k_index[15823] = 74118;
mem_k_index[15824] = 74120;
mem_k_index[15825] = 74123;
mem_k_index[15826] = 74125;
mem_k_index[15827] = 74128;
mem_k_index[15828] = 74130;
mem_k_index[15829] = 74133;
mem_k_index[15830] = 74136;
mem_k_index[15831] = 74138;
mem_k_index[15832] = 74141;
mem_k_index[15833] = 74143;
mem_k_index[15834] = 74146;
mem_k_index[15835] = 74148;
mem_k_index[15836] = 74151;
mem_k_index[15837] = 74153;
mem_k_index[15838] = 74156;
mem_k_index[15839] = 74158;
mem_k_index[15840] = 74161;
mem_k_index[15841] = 74163;
mem_k_index[15842] = 74166;
mem_k_index[15843] = 74168;
mem_k_index[15844] = 74171;
mem_k_index[15845] = 74173;
mem_k_index[15846] = 74176;
mem_k_index[15847] = 74178;
mem_k_index[15848] = 74181;
mem_k_index[15849] = 74183;
mem_k_index[15850] = 74186;
mem_k_index[15851] = 74188;
mem_k_index[15852] = 74191;
mem_k_index[15853] = 74193;
mem_k_index[15854] = 74196;
mem_k_index[15855] = 74198;
mem_k_index[15856] = 74201;
mem_k_index[15857] = 74203;
mem_k_index[15858] = 74206;
mem_k_index[15859] = 74208;
mem_k_index[15860] = 74211;
mem_k_index[15861] = 74213;
mem_k_index[15862] = 74216;
mem_k_index[15863] = 74218;
mem_k_index[15864] = 74221;
mem_k_index[15865] = 74223;
mem_k_index[15866] = 74226;
mem_k_index[15867] = 74228;
mem_k_index[15868] = 74231;
mem_k_index[15869] = 74233;
mem_k_index[15870] = 74236;
mem_k_index[15871] = 74238;
mem_k_index[15872] = 74560;
mem_k_index[15873] = 74562;
mem_k_index[15874] = 74565;
mem_k_index[15875] = 74567;
mem_k_index[15876] = 74570;
mem_k_index[15877] = 74572;
mem_k_index[15878] = 74575;
mem_k_index[15879] = 74577;
mem_k_index[15880] = 74580;
mem_k_index[15881] = 74582;
mem_k_index[15882] = 74585;
mem_k_index[15883] = 74587;
mem_k_index[15884] = 74590;
mem_k_index[15885] = 74592;
mem_k_index[15886] = 74595;
mem_k_index[15887] = 74597;
mem_k_index[15888] = 74600;
mem_k_index[15889] = 74602;
mem_k_index[15890] = 74605;
mem_k_index[15891] = 74607;
mem_k_index[15892] = 74610;
mem_k_index[15893] = 74612;
mem_k_index[15894] = 74615;
mem_k_index[15895] = 74617;
mem_k_index[15896] = 74620;
mem_k_index[15897] = 74622;
mem_k_index[15898] = 74625;
mem_k_index[15899] = 74627;
mem_k_index[15900] = 74630;
mem_k_index[15901] = 74632;
mem_k_index[15902] = 74635;
mem_k_index[15903] = 74637;
mem_k_index[15904] = 74640;
mem_k_index[15905] = 74642;
mem_k_index[15906] = 74645;
mem_k_index[15907] = 74647;
mem_k_index[15908] = 74650;
mem_k_index[15909] = 74652;
mem_k_index[15910] = 74655;
mem_k_index[15911] = 74657;
mem_k_index[15912] = 74660;
mem_k_index[15913] = 74662;
mem_k_index[15914] = 74665;
mem_k_index[15915] = 74668;
mem_k_index[15916] = 74670;
mem_k_index[15917] = 74673;
mem_k_index[15918] = 74675;
mem_k_index[15919] = 74678;
mem_k_index[15920] = 74680;
mem_k_index[15921] = 74683;
mem_k_index[15922] = 74685;
mem_k_index[15923] = 74688;
mem_k_index[15924] = 74690;
mem_k_index[15925] = 74693;
mem_k_index[15926] = 74695;
mem_k_index[15927] = 74698;
mem_k_index[15928] = 74700;
mem_k_index[15929] = 74703;
mem_k_index[15930] = 74705;
mem_k_index[15931] = 74708;
mem_k_index[15932] = 74710;
mem_k_index[15933] = 74713;
mem_k_index[15934] = 74715;
mem_k_index[15935] = 74718;
mem_k_index[15936] = 74720;
mem_k_index[15937] = 74723;
mem_k_index[15938] = 74725;
mem_k_index[15939] = 74728;
mem_k_index[15940] = 74730;
mem_k_index[15941] = 74733;
mem_k_index[15942] = 74735;
mem_k_index[15943] = 74738;
mem_k_index[15944] = 74740;
mem_k_index[15945] = 74743;
mem_k_index[15946] = 74745;
mem_k_index[15947] = 74748;
mem_k_index[15948] = 74750;
mem_k_index[15949] = 74753;
mem_k_index[15950] = 74755;
mem_k_index[15951] = 74758;
mem_k_index[15952] = 74760;
mem_k_index[15953] = 74763;
mem_k_index[15954] = 74765;
mem_k_index[15955] = 74768;
mem_k_index[15956] = 74770;
mem_k_index[15957] = 74773;
mem_k_index[15958] = 74776;
mem_k_index[15959] = 74778;
mem_k_index[15960] = 74781;
mem_k_index[15961] = 74783;
mem_k_index[15962] = 74786;
mem_k_index[15963] = 74788;
mem_k_index[15964] = 74791;
mem_k_index[15965] = 74793;
mem_k_index[15966] = 74796;
mem_k_index[15967] = 74798;
mem_k_index[15968] = 74801;
mem_k_index[15969] = 74803;
mem_k_index[15970] = 74806;
mem_k_index[15971] = 74808;
mem_k_index[15972] = 74811;
mem_k_index[15973] = 74813;
mem_k_index[15974] = 74816;
mem_k_index[15975] = 74818;
mem_k_index[15976] = 74821;
mem_k_index[15977] = 74823;
mem_k_index[15978] = 74826;
mem_k_index[15979] = 74828;
mem_k_index[15980] = 74831;
mem_k_index[15981] = 74833;
mem_k_index[15982] = 74836;
mem_k_index[15983] = 74838;
mem_k_index[15984] = 74841;
mem_k_index[15985] = 74843;
mem_k_index[15986] = 74846;
mem_k_index[15987] = 74848;
mem_k_index[15988] = 74851;
mem_k_index[15989] = 74853;
mem_k_index[15990] = 74856;
mem_k_index[15991] = 74858;
mem_k_index[15992] = 74861;
mem_k_index[15993] = 74863;
mem_k_index[15994] = 74866;
mem_k_index[15995] = 74868;
mem_k_index[15996] = 74871;
mem_k_index[15997] = 74873;
mem_k_index[15998] = 74876;
mem_k_index[15999] = 74878;
mem_k_index[16000] = 75200;
mem_k_index[16001] = 75202;
mem_k_index[16002] = 75205;
mem_k_index[16003] = 75207;
mem_k_index[16004] = 75210;
mem_k_index[16005] = 75212;
mem_k_index[16006] = 75215;
mem_k_index[16007] = 75217;
mem_k_index[16008] = 75220;
mem_k_index[16009] = 75222;
mem_k_index[16010] = 75225;
mem_k_index[16011] = 75227;
mem_k_index[16012] = 75230;
mem_k_index[16013] = 75232;
mem_k_index[16014] = 75235;
mem_k_index[16015] = 75237;
mem_k_index[16016] = 75240;
mem_k_index[16017] = 75242;
mem_k_index[16018] = 75245;
mem_k_index[16019] = 75247;
mem_k_index[16020] = 75250;
mem_k_index[16021] = 75252;
mem_k_index[16022] = 75255;
mem_k_index[16023] = 75257;
mem_k_index[16024] = 75260;
mem_k_index[16025] = 75262;
mem_k_index[16026] = 75265;
mem_k_index[16027] = 75267;
mem_k_index[16028] = 75270;
mem_k_index[16029] = 75272;
mem_k_index[16030] = 75275;
mem_k_index[16031] = 75277;
mem_k_index[16032] = 75280;
mem_k_index[16033] = 75282;
mem_k_index[16034] = 75285;
mem_k_index[16035] = 75287;
mem_k_index[16036] = 75290;
mem_k_index[16037] = 75292;
mem_k_index[16038] = 75295;
mem_k_index[16039] = 75297;
mem_k_index[16040] = 75300;
mem_k_index[16041] = 75302;
mem_k_index[16042] = 75305;
mem_k_index[16043] = 75308;
mem_k_index[16044] = 75310;
mem_k_index[16045] = 75313;
mem_k_index[16046] = 75315;
mem_k_index[16047] = 75318;
mem_k_index[16048] = 75320;
mem_k_index[16049] = 75323;
mem_k_index[16050] = 75325;
mem_k_index[16051] = 75328;
mem_k_index[16052] = 75330;
mem_k_index[16053] = 75333;
mem_k_index[16054] = 75335;
mem_k_index[16055] = 75338;
mem_k_index[16056] = 75340;
mem_k_index[16057] = 75343;
mem_k_index[16058] = 75345;
mem_k_index[16059] = 75348;
mem_k_index[16060] = 75350;
mem_k_index[16061] = 75353;
mem_k_index[16062] = 75355;
mem_k_index[16063] = 75358;
mem_k_index[16064] = 75360;
mem_k_index[16065] = 75363;
mem_k_index[16066] = 75365;
mem_k_index[16067] = 75368;
mem_k_index[16068] = 75370;
mem_k_index[16069] = 75373;
mem_k_index[16070] = 75375;
mem_k_index[16071] = 75378;
mem_k_index[16072] = 75380;
mem_k_index[16073] = 75383;
mem_k_index[16074] = 75385;
mem_k_index[16075] = 75388;
mem_k_index[16076] = 75390;
mem_k_index[16077] = 75393;
mem_k_index[16078] = 75395;
mem_k_index[16079] = 75398;
mem_k_index[16080] = 75400;
mem_k_index[16081] = 75403;
mem_k_index[16082] = 75405;
mem_k_index[16083] = 75408;
mem_k_index[16084] = 75410;
mem_k_index[16085] = 75413;
mem_k_index[16086] = 75416;
mem_k_index[16087] = 75418;
mem_k_index[16088] = 75421;
mem_k_index[16089] = 75423;
mem_k_index[16090] = 75426;
mem_k_index[16091] = 75428;
mem_k_index[16092] = 75431;
mem_k_index[16093] = 75433;
mem_k_index[16094] = 75436;
mem_k_index[16095] = 75438;
mem_k_index[16096] = 75441;
mem_k_index[16097] = 75443;
mem_k_index[16098] = 75446;
mem_k_index[16099] = 75448;
mem_k_index[16100] = 75451;
mem_k_index[16101] = 75453;
mem_k_index[16102] = 75456;
mem_k_index[16103] = 75458;
mem_k_index[16104] = 75461;
mem_k_index[16105] = 75463;
mem_k_index[16106] = 75466;
mem_k_index[16107] = 75468;
mem_k_index[16108] = 75471;
mem_k_index[16109] = 75473;
mem_k_index[16110] = 75476;
mem_k_index[16111] = 75478;
mem_k_index[16112] = 75481;
mem_k_index[16113] = 75483;
mem_k_index[16114] = 75486;
mem_k_index[16115] = 75488;
mem_k_index[16116] = 75491;
mem_k_index[16117] = 75493;
mem_k_index[16118] = 75496;
mem_k_index[16119] = 75498;
mem_k_index[16120] = 75501;
mem_k_index[16121] = 75503;
mem_k_index[16122] = 75506;
mem_k_index[16123] = 75508;
mem_k_index[16124] = 75511;
mem_k_index[16125] = 75513;
mem_k_index[16126] = 75516;
mem_k_index[16127] = 75518;
mem_k_index[16128] = 75840;
mem_k_index[16129] = 75842;
mem_k_index[16130] = 75845;
mem_k_index[16131] = 75847;
mem_k_index[16132] = 75850;
mem_k_index[16133] = 75852;
mem_k_index[16134] = 75855;
mem_k_index[16135] = 75857;
mem_k_index[16136] = 75860;
mem_k_index[16137] = 75862;
mem_k_index[16138] = 75865;
mem_k_index[16139] = 75867;
mem_k_index[16140] = 75870;
mem_k_index[16141] = 75872;
mem_k_index[16142] = 75875;
mem_k_index[16143] = 75877;
mem_k_index[16144] = 75880;
mem_k_index[16145] = 75882;
mem_k_index[16146] = 75885;
mem_k_index[16147] = 75887;
mem_k_index[16148] = 75890;
mem_k_index[16149] = 75892;
mem_k_index[16150] = 75895;
mem_k_index[16151] = 75897;
mem_k_index[16152] = 75900;
mem_k_index[16153] = 75902;
mem_k_index[16154] = 75905;
mem_k_index[16155] = 75907;
mem_k_index[16156] = 75910;
mem_k_index[16157] = 75912;
mem_k_index[16158] = 75915;
mem_k_index[16159] = 75917;
mem_k_index[16160] = 75920;
mem_k_index[16161] = 75922;
mem_k_index[16162] = 75925;
mem_k_index[16163] = 75927;
mem_k_index[16164] = 75930;
mem_k_index[16165] = 75932;
mem_k_index[16166] = 75935;
mem_k_index[16167] = 75937;
mem_k_index[16168] = 75940;
mem_k_index[16169] = 75942;
mem_k_index[16170] = 75945;
mem_k_index[16171] = 75948;
mem_k_index[16172] = 75950;
mem_k_index[16173] = 75953;
mem_k_index[16174] = 75955;
mem_k_index[16175] = 75958;
mem_k_index[16176] = 75960;
mem_k_index[16177] = 75963;
mem_k_index[16178] = 75965;
mem_k_index[16179] = 75968;
mem_k_index[16180] = 75970;
mem_k_index[16181] = 75973;
mem_k_index[16182] = 75975;
mem_k_index[16183] = 75978;
mem_k_index[16184] = 75980;
mem_k_index[16185] = 75983;
mem_k_index[16186] = 75985;
mem_k_index[16187] = 75988;
mem_k_index[16188] = 75990;
mem_k_index[16189] = 75993;
mem_k_index[16190] = 75995;
mem_k_index[16191] = 75998;
mem_k_index[16192] = 76000;
mem_k_index[16193] = 76003;
mem_k_index[16194] = 76005;
mem_k_index[16195] = 76008;
mem_k_index[16196] = 76010;
mem_k_index[16197] = 76013;
mem_k_index[16198] = 76015;
mem_k_index[16199] = 76018;
mem_k_index[16200] = 76020;
mem_k_index[16201] = 76023;
mem_k_index[16202] = 76025;
mem_k_index[16203] = 76028;
mem_k_index[16204] = 76030;
mem_k_index[16205] = 76033;
mem_k_index[16206] = 76035;
mem_k_index[16207] = 76038;
mem_k_index[16208] = 76040;
mem_k_index[16209] = 76043;
mem_k_index[16210] = 76045;
mem_k_index[16211] = 76048;
mem_k_index[16212] = 76050;
mem_k_index[16213] = 76053;
mem_k_index[16214] = 76056;
mem_k_index[16215] = 76058;
mem_k_index[16216] = 76061;
mem_k_index[16217] = 76063;
mem_k_index[16218] = 76066;
mem_k_index[16219] = 76068;
mem_k_index[16220] = 76071;
mem_k_index[16221] = 76073;
mem_k_index[16222] = 76076;
mem_k_index[16223] = 76078;
mem_k_index[16224] = 76081;
mem_k_index[16225] = 76083;
mem_k_index[16226] = 76086;
mem_k_index[16227] = 76088;
mem_k_index[16228] = 76091;
mem_k_index[16229] = 76093;
mem_k_index[16230] = 76096;
mem_k_index[16231] = 76098;
mem_k_index[16232] = 76101;
mem_k_index[16233] = 76103;
mem_k_index[16234] = 76106;
mem_k_index[16235] = 76108;
mem_k_index[16236] = 76111;
mem_k_index[16237] = 76113;
mem_k_index[16238] = 76116;
mem_k_index[16239] = 76118;
mem_k_index[16240] = 76121;
mem_k_index[16241] = 76123;
mem_k_index[16242] = 76126;
mem_k_index[16243] = 76128;
mem_k_index[16244] = 76131;
mem_k_index[16245] = 76133;
mem_k_index[16246] = 76136;
mem_k_index[16247] = 76138;
mem_k_index[16248] = 76141;
mem_k_index[16249] = 76143;
mem_k_index[16250] = 76146;
mem_k_index[16251] = 76148;
mem_k_index[16252] = 76151;
mem_k_index[16253] = 76153;
mem_k_index[16254] = 76156;
mem_k_index[16255] = 76158;
mem_k_index[16256] = 76160;
mem_k_index[16257] = 76162;
mem_k_index[16258] = 76165;
mem_k_index[16259] = 76167;
mem_k_index[16260] = 76170;
mem_k_index[16261] = 76172;
mem_k_index[16262] = 76175;
mem_k_index[16263] = 76177;
mem_k_index[16264] = 76180;
mem_k_index[16265] = 76182;
mem_k_index[16266] = 76185;
mem_k_index[16267] = 76187;
mem_k_index[16268] = 76190;
mem_k_index[16269] = 76192;
mem_k_index[16270] = 76195;
mem_k_index[16271] = 76197;
mem_k_index[16272] = 76200;
mem_k_index[16273] = 76202;
mem_k_index[16274] = 76205;
mem_k_index[16275] = 76207;
mem_k_index[16276] = 76210;
mem_k_index[16277] = 76212;
mem_k_index[16278] = 76215;
mem_k_index[16279] = 76217;
mem_k_index[16280] = 76220;
mem_k_index[16281] = 76222;
mem_k_index[16282] = 76225;
mem_k_index[16283] = 76227;
mem_k_index[16284] = 76230;
mem_k_index[16285] = 76232;
mem_k_index[16286] = 76235;
mem_k_index[16287] = 76237;
mem_k_index[16288] = 76240;
mem_k_index[16289] = 76242;
mem_k_index[16290] = 76245;
mem_k_index[16291] = 76247;
mem_k_index[16292] = 76250;
mem_k_index[16293] = 76252;
mem_k_index[16294] = 76255;
mem_k_index[16295] = 76257;
mem_k_index[16296] = 76260;
mem_k_index[16297] = 76262;
mem_k_index[16298] = 76265;
mem_k_index[16299] = 76268;
mem_k_index[16300] = 76270;
mem_k_index[16301] = 76273;
mem_k_index[16302] = 76275;
mem_k_index[16303] = 76278;
mem_k_index[16304] = 76280;
mem_k_index[16305] = 76283;
mem_k_index[16306] = 76285;
mem_k_index[16307] = 76288;
mem_k_index[16308] = 76290;
mem_k_index[16309] = 76293;
mem_k_index[16310] = 76295;
mem_k_index[16311] = 76298;
mem_k_index[16312] = 76300;
mem_k_index[16313] = 76303;
mem_k_index[16314] = 76305;
mem_k_index[16315] = 76308;
mem_k_index[16316] = 76310;
mem_k_index[16317] = 76313;
mem_k_index[16318] = 76315;
mem_k_index[16319] = 76318;
mem_k_index[16320] = 76320;
mem_k_index[16321] = 76323;
mem_k_index[16322] = 76325;
mem_k_index[16323] = 76328;
mem_k_index[16324] = 76330;
mem_k_index[16325] = 76333;
mem_k_index[16326] = 76335;
mem_k_index[16327] = 76338;
mem_k_index[16328] = 76340;
mem_k_index[16329] = 76343;
mem_k_index[16330] = 76345;
mem_k_index[16331] = 76348;
mem_k_index[16332] = 76350;
mem_k_index[16333] = 76353;
mem_k_index[16334] = 76355;
mem_k_index[16335] = 76358;
mem_k_index[16336] = 76360;
mem_k_index[16337] = 76363;
mem_k_index[16338] = 76365;
mem_k_index[16339] = 76368;
mem_k_index[16340] = 76370;
mem_k_index[16341] = 76373;
mem_k_index[16342] = 76376;
mem_k_index[16343] = 76378;
mem_k_index[16344] = 76381;
mem_k_index[16345] = 76383;
mem_k_index[16346] = 76386;
mem_k_index[16347] = 76388;
mem_k_index[16348] = 76391;
mem_k_index[16349] = 76393;
mem_k_index[16350] = 76396;
mem_k_index[16351] = 76398;
mem_k_index[16352] = 76401;
mem_k_index[16353] = 76403;
mem_k_index[16354] = 76406;
mem_k_index[16355] = 76408;
mem_k_index[16356] = 76411;
mem_k_index[16357] = 76413;
mem_k_index[16358] = 76416;
mem_k_index[16359] = 76418;
mem_k_index[16360] = 76421;
mem_k_index[16361] = 76423;
mem_k_index[16362] = 76426;
mem_k_index[16363] = 76428;
mem_k_index[16364] = 76431;
mem_k_index[16365] = 76433;
mem_k_index[16366] = 76436;
mem_k_index[16367] = 76438;
mem_k_index[16368] = 76441;
mem_k_index[16369] = 76443;
mem_k_index[16370] = 76446;
mem_k_index[16371] = 76448;
mem_k_index[16372] = 76451;
mem_k_index[16373] = 76453;
mem_k_index[16374] = 76456;
mem_k_index[16375] = 76458;
mem_k_index[16376] = 76461;
mem_k_index[16377] = 76463;
mem_k_index[16378] = 76466;
mem_k_index[16379] = 76468;
mem_k_index[16380] = 76471;
mem_k_index[16381] = 76473;
mem_k_index[16382] = 76476;
mem_k_index[16383] = 76478;
end
initial
begin
razn_h_mem[0] = 0;
razn_h_mem[1] = 130;
razn_h_mem[2] = 6;
razn_h_mem[3] = 136;
razn_h_mem[4] = 12;
razn_h_mem[5] = 142;
razn_h_mem[6] = 18;
razn_h_mem[7] = 148;
razn_h_mem[8] = 24;
razn_h_mem[9] = 154;
razn_h_mem[10] = 30;
razn_h_mem[11] = 160;
razn_h_mem[12] = 36;
razn_h_mem[13] = 166;
razn_h_mem[14] = 42;
razn_h_mem[15] = 172;
razn_h_mem[16] = 48;
razn_h_mem[17] = 178;
razn_h_mem[18] = 54;
razn_h_mem[19] = 184;
razn_h_mem[20] = 60;
razn_h_mem[21] = 190;
razn_h_mem[22] = 66;
razn_h_mem[23] = 196;
razn_h_mem[24] = 72;
razn_h_mem[25] = 202;
razn_h_mem[26] = 78;
razn_h_mem[27] = 208;
razn_h_mem[28] = 84;
razn_h_mem[29] = 214;
razn_h_mem[30] = 90;
razn_h_mem[31] = 220;
razn_h_mem[32] = 96;
razn_h_mem[33] = 226;
razn_h_mem[34] = 102;
razn_h_mem[35] = 232;
razn_h_mem[36] = 108;
razn_h_mem[37] = 238;
razn_h_mem[38] = 114;
razn_h_mem[39] = 244;
razn_h_mem[40] = 120;
razn_h_mem[41] = 250;
razn_h_mem[42] = 126;
razn_h_mem[43] = 2;
razn_h_mem[44] = 132;
razn_h_mem[45] = 8;
razn_h_mem[46] = 138;
razn_h_mem[47] = 14;
razn_h_mem[48] = 144;
razn_h_mem[49] = 20;
razn_h_mem[50] = 150;
razn_h_mem[51] = 26;
razn_h_mem[52] = 156;
razn_h_mem[53] = 32;
razn_h_mem[54] = 162;
razn_h_mem[55] = 38;
razn_h_mem[56] = 168;
razn_h_mem[57] = 44;
razn_h_mem[58] = 174;
razn_h_mem[59] = 50;
razn_h_mem[60] = 180;
razn_h_mem[61] = 56;
razn_h_mem[62] = 186;
razn_h_mem[63] = 62;
razn_h_mem[64] = 192;
razn_h_mem[65] = 68;
razn_h_mem[66] = 198;
razn_h_mem[67] = 74;
razn_h_mem[68] = 204;
razn_h_mem[69] = 80;
razn_h_mem[70] = 210;
razn_h_mem[71] = 86;
razn_h_mem[72] = 216;
razn_h_mem[73] = 92;
razn_h_mem[74] = 222;
razn_h_mem[75] = 98;
razn_h_mem[76] = 228;
razn_h_mem[77] = 104;
razn_h_mem[78] = 234;
razn_h_mem[79] = 110;
razn_h_mem[80] = 240;
razn_h_mem[81] = 116;
razn_h_mem[82] = 246;
razn_h_mem[83] = 122;
razn_h_mem[84] = 252;
razn_h_mem[85] = 128;
razn_h_mem[86] = 4;
razn_h_mem[87] = 134;
razn_h_mem[88] = 10;
razn_h_mem[89] = 140;
razn_h_mem[90] = 16;
razn_h_mem[91] = 146;
razn_h_mem[92] = 22;
razn_h_mem[93] = 152;
razn_h_mem[94] = 28;
razn_h_mem[95] = 158;
razn_h_mem[96] = 34;
razn_h_mem[97] = 164;
razn_h_mem[98] = 40;
razn_h_mem[99] = 170;
razn_h_mem[100] = 46;
razn_h_mem[101] = 176;
razn_h_mem[102] = 52;
razn_h_mem[103] = 182;
razn_h_mem[104] = 58;
razn_h_mem[105] = 188;
razn_h_mem[106] = 64;
razn_h_mem[107] = 194;
razn_h_mem[108] = 70;
razn_h_mem[109] = 200;
razn_h_mem[110] = 76;
razn_h_mem[111] = 206;
razn_h_mem[112] = 82;
razn_h_mem[113] = 212;
razn_h_mem[114] = 88;
razn_h_mem[115] = 218;
razn_h_mem[116] = 94;
razn_h_mem[117] = 224;
razn_h_mem[118] = 100;
razn_h_mem[119] = 230;
razn_h_mem[120] = 106;
razn_h_mem[121] = 236;
razn_h_mem[122] = 112;
razn_h_mem[123] = 242;
razn_h_mem[124] = 118;
razn_h_mem[125] = 248;
razn_h_mem[126] = 124;
razn_h_mem[127] = 255;
razn_h_mem[128] = 0;
razn_h_mem[129] = 130;
razn_h_mem[130] = 6;
razn_h_mem[131] = 136;
razn_h_mem[132] = 12;
razn_h_mem[133] = 142;
razn_h_mem[134] = 18;
razn_h_mem[135] = 148;
razn_h_mem[136] = 24;
razn_h_mem[137] = 154;
razn_h_mem[138] = 30;
razn_h_mem[139] = 160;
razn_h_mem[140] = 36;
razn_h_mem[141] = 166;
razn_h_mem[142] = 42;
razn_h_mem[143] = 172;
razn_h_mem[144] = 48;
razn_h_mem[145] = 178;
razn_h_mem[146] = 54;
razn_h_mem[147] = 184;
razn_h_mem[148] = 60;
razn_h_mem[149] = 190;
razn_h_mem[150] = 66;
razn_h_mem[151] = 196;
razn_h_mem[152] = 72;
razn_h_mem[153] = 202;
razn_h_mem[154] = 78;
razn_h_mem[155] = 208;
razn_h_mem[156] = 84;
razn_h_mem[157] = 214;
razn_h_mem[158] = 90;
razn_h_mem[159] = 220;
razn_h_mem[160] = 96;
razn_h_mem[161] = 226;
razn_h_mem[162] = 102;
razn_h_mem[163] = 232;
razn_h_mem[164] = 108;
razn_h_mem[165] = 238;
razn_h_mem[166] = 114;
razn_h_mem[167] = 244;
razn_h_mem[168] = 120;
razn_h_mem[169] = 250;
razn_h_mem[170] = 126;
razn_h_mem[171] = 2;
razn_h_mem[172] = 132;
razn_h_mem[173] = 8;
razn_h_mem[174] = 138;
razn_h_mem[175] = 14;
razn_h_mem[176] = 144;
razn_h_mem[177] = 20;
razn_h_mem[178] = 150;
razn_h_mem[179] = 26;
razn_h_mem[180] = 156;
razn_h_mem[181] = 32;
razn_h_mem[182] = 162;
razn_h_mem[183] = 38;
razn_h_mem[184] = 168;
razn_h_mem[185] = 44;
razn_h_mem[186] = 174;
razn_h_mem[187] = 50;
razn_h_mem[188] = 180;
razn_h_mem[189] = 56;
razn_h_mem[190] = 186;
razn_h_mem[191] = 62;
razn_h_mem[192] = 192;
razn_h_mem[193] = 68;
razn_h_mem[194] = 198;
razn_h_mem[195] = 74;
razn_h_mem[196] = 204;
razn_h_mem[197] = 80;
razn_h_mem[198] = 210;
razn_h_mem[199] = 86;
razn_h_mem[200] = 216;
razn_h_mem[201] = 92;
razn_h_mem[202] = 222;
razn_h_mem[203] = 98;
razn_h_mem[204] = 228;
razn_h_mem[205] = 104;
razn_h_mem[206] = 234;
razn_h_mem[207] = 110;
razn_h_mem[208] = 240;
razn_h_mem[209] = 116;
razn_h_mem[210] = 246;
razn_h_mem[211] = 122;
razn_h_mem[212] = 252;
razn_h_mem[213] = 128;
razn_h_mem[214] = 4;
razn_h_mem[215] = 134;
razn_h_mem[216] = 10;
razn_h_mem[217] = 140;
razn_h_mem[218] = 16;
razn_h_mem[219] = 146;
razn_h_mem[220] = 22;
razn_h_mem[221] = 152;
razn_h_mem[222] = 28;
razn_h_mem[223] = 158;
razn_h_mem[224] = 34;
razn_h_mem[225] = 164;
razn_h_mem[226] = 40;
razn_h_mem[227] = 170;
razn_h_mem[228] = 46;
razn_h_mem[229] = 176;
razn_h_mem[230] = 52;
razn_h_mem[231] = 182;
razn_h_mem[232] = 58;
razn_h_mem[233] = 188;
razn_h_mem[234] = 64;
razn_h_mem[235] = 194;
razn_h_mem[236] = 70;
razn_h_mem[237] = 200;
razn_h_mem[238] = 76;
razn_h_mem[239] = 206;
razn_h_mem[240] = 82;
razn_h_mem[241] = 212;
razn_h_mem[242] = 88;
razn_h_mem[243] = 218;
razn_h_mem[244] = 94;
razn_h_mem[245] = 224;
razn_h_mem[246] = 100;
razn_h_mem[247] = 230;
razn_h_mem[248] = 106;
razn_h_mem[249] = 236;
razn_h_mem[250] = 112;
razn_h_mem[251] = 242;
razn_h_mem[252] = 118;
razn_h_mem[253] = 248;
razn_h_mem[254] = 124;
razn_h_mem[255] = 255;
razn_h_mem[256] = 0;
razn_h_mem[257] = 130;
razn_h_mem[258] = 6;
razn_h_mem[259] = 136;
razn_h_mem[260] = 12;
razn_h_mem[261] = 142;
razn_h_mem[262] = 18;
razn_h_mem[263] = 148;
razn_h_mem[264] = 24;
razn_h_mem[265] = 154;
razn_h_mem[266] = 30;
razn_h_mem[267] = 160;
razn_h_mem[268] = 36;
razn_h_mem[269] = 166;
razn_h_mem[270] = 42;
razn_h_mem[271] = 172;
razn_h_mem[272] = 48;
razn_h_mem[273] = 178;
razn_h_mem[274] = 54;
razn_h_mem[275] = 184;
razn_h_mem[276] = 60;
razn_h_mem[277] = 190;
razn_h_mem[278] = 66;
razn_h_mem[279] = 196;
razn_h_mem[280] = 72;
razn_h_mem[281] = 202;
razn_h_mem[282] = 78;
razn_h_mem[283] = 208;
razn_h_mem[284] = 84;
razn_h_mem[285] = 214;
razn_h_mem[286] = 90;
razn_h_mem[287] = 220;
razn_h_mem[288] = 96;
razn_h_mem[289] = 226;
razn_h_mem[290] = 102;
razn_h_mem[291] = 232;
razn_h_mem[292] = 108;
razn_h_mem[293] = 238;
razn_h_mem[294] = 114;
razn_h_mem[295] = 244;
razn_h_mem[296] = 120;
razn_h_mem[297] = 250;
razn_h_mem[298] = 126;
razn_h_mem[299] = 2;
razn_h_mem[300] = 132;
razn_h_mem[301] = 8;
razn_h_mem[302] = 138;
razn_h_mem[303] = 14;
razn_h_mem[304] = 144;
razn_h_mem[305] = 20;
razn_h_mem[306] = 150;
razn_h_mem[307] = 26;
razn_h_mem[308] = 156;
razn_h_mem[309] = 32;
razn_h_mem[310] = 162;
razn_h_mem[311] = 38;
razn_h_mem[312] = 168;
razn_h_mem[313] = 44;
razn_h_mem[314] = 174;
razn_h_mem[315] = 50;
razn_h_mem[316] = 180;
razn_h_mem[317] = 56;
razn_h_mem[318] = 186;
razn_h_mem[319] = 62;
razn_h_mem[320] = 192;
razn_h_mem[321] = 68;
razn_h_mem[322] = 198;
razn_h_mem[323] = 74;
razn_h_mem[324] = 204;
razn_h_mem[325] = 80;
razn_h_mem[326] = 210;
razn_h_mem[327] = 86;
razn_h_mem[328] = 216;
razn_h_mem[329] = 92;
razn_h_mem[330] = 222;
razn_h_mem[331] = 98;
razn_h_mem[332] = 228;
razn_h_mem[333] = 104;
razn_h_mem[334] = 234;
razn_h_mem[335] = 110;
razn_h_mem[336] = 240;
razn_h_mem[337] = 116;
razn_h_mem[338] = 246;
razn_h_mem[339] = 122;
razn_h_mem[340] = 252;
razn_h_mem[341] = 128;
razn_h_mem[342] = 4;
razn_h_mem[343] = 134;
razn_h_mem[344] = 10;
razn_h_mem[345] = 140;
razn_h_mem[346] = 16;
razn_h_mem[347] = 146;
razn_h_mem[348] = 22;
razn_h_mem[349] = 152;
razn_h_mem[350] = 28;
razn_h_mem[351] = 158;
razn_h_mem[352] = 34;
razn_h_mem[353] = 164;
razn_h_mem[354] = 40;
razn_h_mem[355] = 170;
razn_h_mem[356] = 46;
razn_h_mem[357] = 176;
razn_h_mem[358] = 52;
razn_h_mem[359] = 182;
razn_h_mem[360] = 58;
razn_h_mem[361] = 188;
razn_h_mem[362] = 64;
razn_h_mem[363] = 194;
razn_h_mem[364] = 70;
razn_h_mem[365] = 200;
razn_h_mem[366] = 76;
razn_h_mem[367] = 206;
razn_h_mem[368] = 82;
razn_h_mem[369] = 212;
razn_h_mem[370] = 88;
razn_h_mem[371] = 218;
razn_h_mem[372] = 94;
razn_h_mem[373] = 224;
razn_h_mem[374] = 100;
razn_h_mem[375] = 230;
razn_h_mem[376] = 106;
razn_h_mem[377] = 236;
razn_h_mem[378] = 112;
razn_h_mem[379] = 242;
razn_h_mem[380] = 118;
razn_h_mem[381] = 248;
razn_h_mem[382] = 124;
razn_h_mem[383] = 255;
razn_h_mem[384] = 0;
razn_h_mem[385] = 130;
razn_h_mem[386] = 6;
razn_h_mem[387] = 136;
razn_h_mem[388] = 12;
razn_h_mem[389] = 142;
razn_h_mem[390] = 18;
razn_h_mem[391] = 148;
razn_h_mem[392] = 24;
razn_h_mem[393] = 154;
razn_h_mem[394] = 30;
razn_h_mem[395] = 160;
razn_h_mem[396] = 36;
razn_h_mem[397] = 166;
razn_h_mem[398] = 42;
razn_h_mem[399] = 172;
razn_h_mem[400] = 48;
razn_h_mem[401] = 178;
razn_h_mem[402] = 54;
razn_h_mem[403] = 184;
razn_h_mem[404] = 60;
razn_h_mem[405] = 190;
razn_h_mem[406] = 66;
razn_h_mem[407] = 196;
razn_h_mem[408] = 72;
razn_h_mem[409] = 202;
razn_h_mem[410] = 78;
razn_h_mem[411] = 208;
razn_h_mem[412] = 84;
razn_h_mem[413] = 214;
razn_h_mem[414] = 90;
razn_h_mem[415] = 220;
razn_h_mem[416] = 96;
razn_h_mem[417] = 226;
razn_h_mem[418] = 102;
razn_h_mem[419] = 232;
razn_h_mem[420] = 108;
razn_h_mem[421] = 238;
razn_h_mem[422] = 114;
razn_h_mem[423] = 244;
razn_h_mem[424] = 120;
razn_h_mem[425] = 250;
razn_h_mem[426] = 126;
razn_h_mem[427] = 2;
razn_h_mem[428] = 132;
razn_h_mem[429] = 8;
razn_h_mem[430] = 138;
razn_h_mem[431] = 14;
razn_h_mem[432] = 144;
razn_h_mem[433] = 20;
razn_h_mem[434] = 150;
razn_h_mem[435] = 26;
razn_h_mem[436] = 156;
razn_h_mem[437] = 32;
razn_h_mem[438] = 162;
razn_h_mem[439] = 38;
razn_h_mem[440] = 168;
razn_h_mem[441] = 44;
razn_h_mem[442] = 174;
razn_h_mem[443] = 50;
razn_h_mem[444] = 180;
razn_h_mem[445] = 56;
razn_h_mem[446] = 186;
razn_h_mem[447] = 62;
razn_h_mem[448] = 192;
razn_h_mem[449] = 68;
razn_h_mem[450] = 198;
razn_h_mem[451] = 74;
razn_h_mem[452] = 204;
razn_h_mem[453] = 80;
razn_h_mem[454] = 210;
razn_h_mem[455] = 86;
razn_h_mem[456] = 216;
razn_h_mem[457] = 92;
razn_h_mem[458] = 222;
razn_h_mem[459] = 98;
razn_h_mem[460] = 228;
razn_h_mem[461] = 104;
razn_h_mem[462] = 234;
razn_h_mem[463] = 110;
razn_h_mem[464] = 240;
razn_h_mem[465] = 116;
razn_h_mem[466] = 246;
razn_h_mem[467] = 122;
razn_h_mem[468] = 252;
razn_h_mem[469] = 128;
razn_h_mem[470] = 4;
razn_h_mem[471] = 134;
razn_h_mem[472] = 10;
razn_h_mem[473] = 140;
razn_h_mem[474] = 16;
razn_h_mem[475] = 146;
razn_h_mem[476] = 22;
razn_h_mem[477] = 152;
razn_h_mem[478] = 28;
razn_h_mem[479] = 158;
razn_h_mem[480] = 34;
razn_h_mem[481] = 164;
razn_h_mem[482] = 40;
razn_h_mem[483] = 170;
razn_h_mem[484] = 46;
razn_h_mem[485] = 176;
razn_h_mem[486] = 52;
razn_h_mem[487] = 182;
razn_h_mem[488] = 58;
razn_h_mem[489] = 188;
razn_h_mem[490] = 64;
razn_h_mem[491] = 194;
razn_h_mem[492] = 70;
razn_h_mem[493] = 200;
razn_h_mem[494] = 76;
razn_h_mem[495] = 206;
razn_h_mem[496] = 82;
razn_h_mem[497] = 212;
razn_h_mem[498] = 88;
razn_h_mem[499] = 218;
razn_h_mem[500] = 94;
razn_h_mem[501] = 224;
razn_h_mem[502] = 100;
razn_h_mem[503] = 230;
razn_h_mem[504] = 106;
razn_h_mem[505] = 236;
razn_h_mem[506] = 112;
razn_h_mem[507] = 242;
razn_h_mem[508] = 118;
razn_h_mem[509] = 248;
razn_h_mem[510] = 124;
razn_h_mem[511] = 255;
razn_h_mem[512] = 0;
razn_h_mem[513] = 130;
razn_h_mem[514] = 6;
razn_h_mem[515] = 136;
razn_h_mem[516] = 12;
razn_h_mem[517] = 142;
razn_h_mem[518] = 18;
razn_h_mem[519] = 148;
razn_h_mem[520] = 24;
razn_h_mem[521] = 154;
razn_h_mem[522] = 30;
razn_h_mem[523] = 160;
razn_h_mem[524] = 36;
razn_h_mem[525] = 166;
razn_h_mem[526] = 42;
razn_h_mem[527] = 172;
razn_h_mem[528] = 48;
razn_h_mem[529] = 178;
razn_h_mem[530] = 54;
razn_h_mem[531] = 184;
razn_h_mem[532] = 60;
razn_h_mem[533] = 190;
razn_h_mem[534] = 66;
razn_h_mem[535] = 196;
razn_h_mem[536] = 72;
razn_h_mem[537] = 202;
razn_h_mem[538] = 78;
razn_h_mem[539] = 208;
razn_h_mem[540] = 84;
razn_h_mem[541] = 214;
razn_h_mem[542] = 90;
razn_h_mem[543] = 220;
razn_h_mem[544] = 96;
razn_h_mem[545] = 226;
razn_h_mem[546] = 102;
razn_h_mem[547] = 232;
razn_h_mem[548] = 108;
razn_h_mem[549] = 238;
razn_h_mem[550] = 114;
razn_h_mem[551] = 244;
razn_h_mem[552] = 120;
razn_h_mem[553] = 250;
razn_h_mem[554] = 126;
razn_h_mem[555] = 2;
razn_h_mem[556] = 132;
razn_h_mem[557] = 8;
razn_h_mem[558] = 138;
razn_h_mem[559] = 14;
razn_h_mem[560] = 144;
razn_h_mem[561] = 20;
razn_h_mem[562] = 150;
razn_h_mem[563] = 26;
razn_h_mem[564] = 156;
razn_h_mem[565] = 32;
razn_h_mem[566] = 162;
razn_h_mem[567] = 38;
razn_h_mem[568] = 168;
razn_h_mem[569] = 44;
razn_h_mem[570] = 174;
razn_h_mem[571] = 50;
razn_h_mem[572] = 180;
razn_h_mem[573] = 56;
razn_h_mem[574] = 186;
razn_h_mem[575] = 62;
razn_h_mem[576] = 192;
razn_h_mem[577] = 68;
razn_h_mem[578] = 198;
razn_h_mem[579] = 74;
razn_h_mem[580] = 204;
razn_h_mem[581] = 80;
razn_h_mem[582] = 210;
razn_h_mem[583] = 86;
razn_h_mem[584] = 216;
razn_h_mem[585] = 92;
razn_h_mem[586] = 222;
razn_h_mem[587] = 98;
razn_h_mem[588] = 228;
razn_h_mem[589] = 104;
razn_h_mem[590] = 234;
razn_h_mem[591] = 110;
razn_h_mem[592] = 240;
razn_h_mem[593] = 116;
razn_h_mem[594] = 246;
razn_h_mem[595] = 122;
razn_h_mem[596] = 252;
razn_h_mem[597] = 128;
razn_h_mem[598] = 4;
razn_h_mem[599] = 134;
razn_h_mem[600] = 10;
razn_h_mem[601] = 140;
razn_h_mem[602] = 16;
razn_h_mem[603] = 146;
razn_h_mem[604] = 22;
razn_h_mem[605] = 152;
razn_h_mem[606] = 28;
razn_h_mem[607] = 158;
razn_h_mem[608] = 34;
razn_h_mem[609] = 164;
razn_h_mem[610] = 40;
razn_h_mem[611] = 170;
razn_h_mem[612] = 46;
razn_h_mem[613] = 176;
razn_h_mem[614] = 52;
razn_h_mem[615] = 182;
razn_h_mem[616] = 58;
razn_h_mem[617] = 188;
razn_h_mem[618] = 64;
razn_h_mem[619] = 194;
razn_h_mem[620] = 70;
razn_h_mem[621] = 200;
razn_h_mem[622] = 76;
razn_h_mem[623] = 206;
razn_h_mem[624] = 82;
razn_h_mem[625] = 212;
razn_h_mem[626] = 88;
razn_h_mem[627] = 218;
razn_h_mem[628] = 94;
razn_h_mem[629] = 224;
razn_h_mem[630] = 100;
razn_h_mem[631] = 230;
razn_h_mem[632] = 106;
razn_h_mem[633] = 236;
razn_h_mem[634] = 112;
razn_h_mem[635] = 242;
razn_h_mem[636] = 118;
razn_h_mem[637] = 248;
razn_h_mem[638] = 124;
razn_h_mem[639] = 255;
razn_h_mem[640] = 0;
razn_h_mem[641] = 130;
razn_h_mem[642] = 6;
razn_h_mem[643] = 136;
razn_h_mem[644] = 12;
razn_h_mem[645] = 142;
razn_h_mem[646] = 18;
razn_h_mem[647] = 148;
razn_h_mem[648] = 24;
razn_h_mem[649] = 154;
razn_h_mem[650] = 30;
razn_h_mem[651] = 160;
razn_h_mem[652] = 36;
razn_h_mem[653] = 166;
razn_h_mem[654] = 42;
razn_h_mem[655] = 172;
razn_h_mem[656] = 48;
razn_h_mem[657] = 178;
razn_h_mem[658] = 54;
razn_h_mem[659] = 184;
razn_h_mem[660] = 60;
razn_h_mem[661] = 190;
razn_h_mem[662] = 66;
razn_h_mem[663] = 196;
razn_h_mem[664] = 72;
razn_h_mem[665] = 202;
razn_h_mem[666] = 78;
razn_h_mem[667] = 208;
razn_h_mem[668] = 84;
razn_h_mem[669] = 214;
razn_h_mem[670] = 90;
razn_h_mem[671] = 220;
razn_h_mem[672] = 96;
razn_h_mem[673] = 226;
razn_h_mem[674] = 102;
razn_h_mem[675] = 232;
razn_h_mem[676] = 108;
razn_h_mem[677] = 238;
razn_h_mem[678] = 114;
razn_h_mem[679] = 244;
razn_h_mem[680] = 120;
razn_h_mem[681] = 250;
razn_h_mem[682] = 126;
razn_h_mem[683] = 2;
razn_h_mem[684] = 132;
razn_h_mem[685] = 8;
razn_h_mem[686] = 138;
razn_h_mem[687] = 14;
razn_h_mem[688] = 144;
razn_h_mem[689] = 20;
razn_h_mem[690] = 150;
razn_h_mem[691] = 26;
razn_h_mem[692] = 156;
razn_h_mem[693] = 32;
razn_h_mem[694] = 162;
razn_h_mem[695] = 38;
razn_h_mem[696] = 168;
razn_h_mem[697] = 44;
razn_h_mem[698] = 174;
razn_h_mem[699] = 50;
razn_h_mem[700] = 180;
razn_h_mem[701] = 56;
razn_h_mem[702] = 186;
razn_h_mem[703] = 62;
razn_h_mem[704] = 192;
razn_h_mem[705] = 68;
razn_h_mem[706] = 198;
razn_h_mem[707] = 74;
razn_h_mem[708] = 204;
razn_h_mem[709] = 80;
razn_h_mem[710] = 210;
razn_h_mem[711] = 86;
razn_h_mem[712] = 216;
razn_h_mem[713] = 92;
razn_h_mem[714] = 222;
razn_h_mem[715] = 98;
razn_h_mem[716] = 228;
razn_h_mem[717] = 104;
razn_h_mem[718] = 234;
razn_h_mem[719] = 110;
razn_h_mem[720] = 240;
razn_h_mem[721] = 116;
razn_h_mem[722] = 246;
razn_h_mem[723] = 122;
razn_h_mem[724] = 252;
razn_h_mem[725] = 128;
razn_h_mem[726] = 4;
razn_h_mem[727] = 134;
razn_h_mem[728] = 10;
razn_h_mem[729] = 140;
razn_h_mem[730] = 16;
razn_h_mem[731] = 146;
razn_h_mem[732] = 22;
razn_h_mem[733] = 152;
razn_h_mem[734] = 28;
razn_h_mem[735] = 158;
razn_h_mem[736] = 34;
razn_h_mem[737] = 164;
razn_h_mem[738] = 40;
razn_h_mem[739] = 170;
razn_h_mem[740] = 46;
razn_h_mem[741] = 176;
razn_h_mem[742] = 52;
razn_h_mem[743] = 182;
razn_h_mem[744] = 58;
razn_h_mem[745] = 188;
razn_h_mem[746] = 64;
razn_h_mem[747] = 194;
razn_h_mem[748] = 70;
razn_h_mem[749] = 200;
razn_h_mem[750] = 76;
razn_h_mem[751] = 206;
razn_h_mem[752] = 82;
razn_h_mem[753] = 212;
razn_h_mem[754] = 88;
razn_h_mem[755] = 218;
razn_h_mem[756] = 94;
razn_h_mem[757] = 224;
razn_h_mem[758] = 100;
razn_h_mem[759] = 230;
razn_h_mem[760] = 106;
razn_h_mem[761] = 236;
razn_h_mem[762] = 112;
razn_h_mem[763] = 242;
razn_h_mem[764] = 118;
razn_h_mem[765] = 248;
razn_h_mem[766] = 124;
razn_h_mem[767] = 255;
razn_h_mem[768] = 0;
razn_h_mem[769] = 130;
razn_h_mem[770] = 6;
razn_h_mem[771] = 136;
razn_h_mem[772] = 12;
razn_h_mem[773] = 142;
razn_h_mem[774] = 18;
razn_h_mem[775] = 148;
razn_h_mem[776] = 24;
razn_h_mem[777] = 154;
razn_h_mem[778] = 30;
razn_h_mem[779] = 160;
razn_h_mem[780] = 36;
razn_h_mem[781] = 166;
razn_h_mem[782] = 42;
razn_h_mem[783] = 172;
razn_h_mem[784] = 48;
razn_h_mem[785] = 178;
razn_h_mem[786] = 54;
razn_h_mem[787] = 184;
razn_h_mem[788] = 60;
razn_h_mem[789] = 190;
razn_h_mem[790] = 66;
razn_h_mem[791] = 196;
razn_h_mem[792] = 72;
razn_h_mem[793] = 202;
razn_h_mem[794] = 78;
razn_h_mem[795] = 208;
razn_h_mem[796] = 84;
razn_h_mem[797] = 214;
razn_h_mem[798] = 90;
razn_h_mem[799] = 220;
razn_h_mem[800] = 96;
razn_h_mem[801] = 226;
razn_h_mem[802] = 102;
razn_h_mem[803] = 232;
razn_h_mem[804] = 108;
razn_h_mem[805] = 238;
razn_h_mem[806] = 114;
razn_h_mem[807] = 244;
razn_h_mem[808] = 120;
razn_h_mem[809] = 250;
razn_h_mem[810] = 126;
razn_h_mem[811] = 2;
razn_h_mem[812] = 132;
razn_h_mem[813] = 8;
razn_h_mem[814] = 138;
razn_h_mem[815] = 14;
razn_h_mem[816] = 144;
razn_h_mem[817] = 20;
razn_h_mem[818] = 150;
razn_h_mem[819] = 26;
razn_h_mem[820] = 156;
razn_h_mem[821] = 32;
razn_h_mem[822] = 162;
razn_h_mem[823] = 38;
razn_h_mem[824] = 168;
razn_h_mem[825] = 44;
razn_h_mem[826] = 174;
razn_h_mem[827] = 50;
razn_h_mem[828] = 180;
razn_h_mem[829] = 56;
razn_h_mem[830] = 186;
razn_h_mem[831] = 62;
razn_h_mem[832] = 192;
razn_h_mem[833] = 68;
razn_h_mem[834] = 198;
razn_h_mem[835] = 74;
razn_h_mem[836] = 204;
razn_h_mem[837] = 80;
razn_h_mem[838] = 210;
razn_h_mem[839] = 86;
razn_h_mem[840] = 216;
razn_h_mem[841] = 92;
razn_h_mem[842] = 222;
razn_h_mem[843] = 98;
razn_h_mem[844] = 228;
razn_h_mem[845] = 104;
razn_h_mem[846] = 234;
razn_h_mem[847] = 110;
razn_h_mem[848] = 240;
razn_h_mem[849] = 116;
razn_h_mem[850] = 246;
razn_h_mem[851] = 122;
razn_h_mem[852] = 252;
razn_h_mem[853] = 128;
razn_h_mem[854] = 4;
razn_h_mem[855] = 134;
razn_h_mem[856] = 10;
razn_h_mem[857] = 140;
razn_h_mem[858] = 16;
razn_h_mem[859] = 146;
razn_h_mem[860] = 22;
razn_h_mem[861] = 152;
razn_h_mem[862] = 28;
razn_h_mem[863] = 158;
razn_h_mem[864] = 34;
razn_h_mem[865] = 164;
razn_h_mem[866] = 40;
razn_h_mem[867] = 170;
razn_h_mem[868] = 46;
razn_h_mem[869] = 176;
razn_h_mem[870] = 52;
razn_h_mem[871] = 182;
razn_h_mem[872] = 58;
razn_h_mem[873] = 188;
razn_h_mem[874] = 64;
razn_h_mem[875] = 194;
razn_h_mem[876] = 70;
razn_h_mem[877] = 200;
razn_h_mem[878] = 76;
razn_h_mem[879] = 206;
razn_h_mem[880] = 82;
razn_h_mem[881] = 212;
razn_h_mem[882] = 88;
razn_h_mem[883] = 218;
razn_h_mem[884] = 94;
razn_h_mem[885] = 224;
razn_h_mem[886] = 100;
razn_h_mem[887] = 230;
razn_h_mem[888] = 106;
razn_h_mem[889] = 236;
razn_h_mem[890] = 112;
razn_h_mem[891] = 242;
razn_h_mem[892] = 118;
razn_h_mem[893] = 248;
razn_h_mem[894] = 124;
razn_h_mem[895] = 255;
razn_h_mem[896] = 0;
razn_h_mem[897] = 130;
razn_h_mem[898] = 6;
razn_h_mem[899] = 136;
razn_h_mem[900] = 12;
razn_h_mem[901] = 142;
razn_h_mem[902] = 18;
razn_h_mem[903] = 148;
razn_h_mem[904] = 24;
razn_h_mem[905] = 154;
razn_h_mem[906] = 30;
razn_h_mem[907] = 160;
razn_h_mem[908] = 36;
razn_h_mem[909] = 166;
razn_h_mem[910] = 42;
razn_h_mem[911] = 172;
razn_h_mem[912] = 48;
razn_h_mem[913] = 178;
razn_h_mem[914] = 54;
razn_h_mem[915] = 184;
razn_h_mem[916] = 60;
razn_h_mem[917] = 190;
razn_h_mem[918] = 66;
razn_h_mem[919] = 196;
razn_h_mem[920] = 72;
razn_h_mem[921] = 202;
razn_h_mem[922] = 78;
razn_h_mem[923] = 208;
razn_h_mem[924] = 84;
razn_h_mem[925] = 214;
razn_h_mem[926] = 90;
razn_h_mem[927] = 220;
razn_h_mem[928] = 96;
razn_h_mem[929] = 226;
razn_h_mem[930] = 102;
razn_h_mem[931] = 232;
razn_h_mem[932] = 108;
razn_h_mem[933] = 238;
razn_h_mem[934] = 114;
razn_h_mem[935] = 244;
razn_h_mem[936] = 120;
razn_h_mem[937] = 250;
razn_h_mem[938] = 126;
razn_h_mem[939] = 2;
razn_h_mem[940] = 132;
razn_h_mem[941] = 8;
razn_h_mem[942] = 138;
razn_h_mem[943] = 14;
razn_h_mem[944] = 144;
razn_h_mem[945] = 20;
razn_h_mem[946] = 150;
razn_h_mem[947] = 26;
razn_h_mem[948] = 156;
razn_h_mem[949] = 32;
razn_h_mem[950] = 162;
razn_h_mem[951] = 38;
razn_h_mem[952] = 168;
razn_h_mem[953] = 44;
razn_h_mem[954] = 174;
razn_h_mem[955] = 50;
razn_h_mem[956] = 180;
razn_h_mem[957] = 56;
razn_h_mem[958] = 186;
razn_h_mem[959] = 62;
razn_h_mem[960] = 192;
razn_h_mem[961] = 68;
razn_h_mem[962] = 198;
razn_h_mem[963] = 74;
razn_h_mem[964] = 204;
razn_h_mem[965] = 80;
razn_h_mem[966] = 210;
razn_h_mem[967] = 86;
razn_h_mem[968] = 216;
razn_h_mem[969] = 92;
razn_h_mem[970] = 222;
razn_h_mem[971] = 98;
razn_h_mem[972] = 228;
razn_h_mem[973] = 104;
razn_h_mem[974] = 234;
razn_h_mem[975] = 110;
razn_h_mem[976] = 240;
razn_h_mem[977] = 116;
razn_h_mem[978] = 246;
razn_h_mem[979] = 122;
razn_h_mem[980] = 252;
razn_h_mem[981] = 128;
razn_h_mem[982] = 4;
razn_h_mem[983] = 134;
razn_h_mem[984] = 10;
razn_h_mem[985] = 140;
razn_h_mem[986] = 16;
razn_h_mem[987] = 146;
razn_h_mem[988] = 22;
razn_h_mem[989] = 152;
razn_h_mem[990] = 28;
razn_h_mem[991] = 158;
razn_h_mem[992] = 34;
razn_h_mem[993] = 164;
razn_h_mem[994] = 40;
razn_h_mem[995] = 170;
razn_h_mem[996] = 46;
razn_h_mem[997] = 176;
razn_h_mem[998] = 52;
razn_h_mem[999] = 182;
razn_h_mem[1000] = 58;
razn_h_mem[1001] = 188;
razn_h_mem[1002] = 64;
razn_h_mem[1003] = 194;
razn_h_mem[1004] = 70;
razn_h_mem[1005] = 200;
razn_h_mem[1006] = 76;
razn_h_mem[1007] = 206;
razn_h_mem[1008] = 82;
razn_h_mem[1009] = 212;
razn_h_mem[1010] = 88;
razn_h_mem[1011] = 218;
razn_h_mem[1012] = 94;
razn_h_mem[1013] = 224;
razn_h_mem[1014] = 100;
razn_h_mem[1015] = 230;
razn_h_mem[1016] = 106;
razn_h_mem[1017] = 236;
razn_h_mem[1018] = 112;
razn_h_mem[1019] = 242;
razn_h_mem[1020] = 118;
razn_h_mem[1021] = 248;
razn_h_mem[1022] = 124;
razn_h_mem[1023] = 255;
razn_h_mem[1024] = 0;
razn_h_mem[1025] = 130;
razn_h_mem[1026] = 6;
razn_h_mem[1027] = 136;
razn_h_mem[1028] = 12;
razn_h_mem[1029] = 142;
razn_h_mem[1030] = 18;
razn_h_mem[1031] = 148;
razn_h_mem[1032] = 24;
razn_h_mem[1033] = 154;
razn_h_mem[1034] = 30;
razn_h_mem[1035] = 160;
razn_h_mem[1036] = 36;
razn_h_mem[1037] = 166;
razn_h_mem[1038] = 42;
razn_h_mem[1039] = 172;
razn_h_mem[1040] = 48;
razn_h_mem[1041] = 178;
razn_h_mem[1042] = 54;
razn_h_mem[1043] = 184;
razn_h_mem[1044] = 60;
razn_h_mem[1045] = 190;
razn_h_mem[1046] = 66;
razn_h_mem[1047] = 196;
razn_h_mem[1048] = 72;
razn_h_mem[1049] = 202;
razn_h_mem[1050] = 78;
razn_h_mem[1051] = 208;
razn_h_mem[1052] = 84;
razn_h_mem[1053] = 214;
razn_h_mem[1054] = 90;
razn_h_mem[1055] = 220;
razn_h_mem[1056] = 96;
razn_h_mem[1057] = 226;
razn_h_mem[1058] = 102;
razn_h_mem[1059] = 232;
razn_h_mem[1060] = 108;
razn_h_mem[1061] = 238;
razn_h_mem[1062] = 114;
razn_h_mem[1063] = 244;
razn_h_mem[1064] = 120;
razn_h_mem[1065] = 250;
razn_h_mem[1066] = 126;
razn_h_mem[1067] = 2;
razn_h_mem[1068] = 132;
razn_h_mem[1069] = 8;
razn_h_mem[1070] = 138;
razn_h_mem[1071] = 14;
razn_h_mem[1072] = 144;
razn_h_mem[1073] = 20;
razn_h_mem[1074] = 150;
razn_h_mem[1075] = 26;
razn_h_mem[1076] = 156;
razn_h_mem[1077] = 32;
razn_h_mem[1078] = 162;
razn_h_mem[1079] = 38;
razn_h_mem[1080] = 168;
razn_h_mem[1081] = 44;
razn_h_mem[1082] = 174;
razn_h_mem[1083] = 50;
razn_h_mem[1084] = 180;
razn_h_mem[1085] = 56;
razn_h_mem[1086] = 186;
razn_h_mem[1087] = 62;
razn_h_mem[1088] = 192;
razn_h_mem[1089] = 68;
razn_h_mem[1090] = 198;
razn_h_mem[1091] = 74;
razn_h_mem[1092] = 204;
razn_h_mem[1093] = 80;
razn_h_mem[1094] = 210;
razn_h_mem[1095] = 86;
razn_h_mem[1096] = 216;
razn_h_mem[1097] = 92;
razn_h_mem[1098] = 222;
razn_h_mem[1099] = 98;
razn_h_mem[1100] = 228;
razn_h_mem[1101] = 104;
razn_h_mem[1102] = 234;
razn_h_mem[1103] = 110;
razn_h_mem[1104] = 240;
razn_h_mem[1105] = 116;
razn_h_mem[1106] = 246;
razn_h_mem[1107] = 122;
razn_h_mem[1108] = 252;
razn_h_mem[1109] = 128;
razn_h_mem[1110] = 4;
razn_h_mem[1111] = 134;
razn_h_mem[1112] = 10;
razn_h_mem[1113] = 140;
razn_h_mem[1114] = 16;
razn_h_mem[1115] = 146;
razn_h_mem[1116] = 22;
razn_h_mem[1117] = 152;
razn_h_mem[1118] = 28;
razn_h_mem[1119] = 158;
razn_h_mem[1120] = 34;
razn_h_mem[1121] = 164;
razn_h_mem[1122] = 40;
razn_h_mem[1123] = 170;
razn_h_mem[1124] = 46;
razn_h_mem[1125] = 176;
razn_h_mem[1126] = 52;
razn_h_mem[1127] = 182;
razn_h_mem[1128] = 58;
razn_h_mem[1129] = 188;
razn_h_mem[1130] = 64;
razn_h_mem[1131] = 194;
razn_h_mem[1132] = 70;
razn_h_mem[1133] = 200;
razn_h_mem[1134] = 76;
razn_h_mem[1135] = 206;
razn_h_mem[1136] = 82;
razn_h_mem[1137] = 212;
razn_h_mem[1138] = 88;
razn_h_mem[1139] = 218;
razn_h_mem[1140] = 94;
razn_h_mem[1141] = 224;
razn_h_mem[1142] = 100;
razn_h_mem[1143] = 230;
razn_h_mem[1144] = 106;
razn_h_mem[1145] = 236;
razn_h_mem[1146] = 112;
razn_h_mem[1147] = 242;
razn_h_mem[1148] = 118;
razn_h_mem[1149] = 248;
razn_h_mem[1150] = 124;
razn_h_mem[1151] = 255;
razn_h_mem[1152] = 0;
razn_h_mem[1153] = 130;
razn_h_mem[1154] = 6;
razn_h_mem[1155] = 136;
razn_h_mem[1156] = 12;
razn_h_mem[1157] = 142;
razn_h_mem[1158] = 18;
razn_h_mem[1159] = 148;
razn_h_mem[1160] = 24;
razn_h_mem[1161] = 154;
razn_h_mem[1162] = 30;
razn_h_mem[1163] = 160;
razn_h_mem[1164] = 36;
razn_h_mem[1165] = 166;
razn_h_mem[1166] = 42;
razn_h_mem[1167] = 172;
razn_h_mem[1168] = 48;
razn_h_mem[1169] = 178;
razn_h_mem[1170] = 54;
razn_h_mem[1171] = 184;
razn_h_mem[1172] = 60;
razn_h_mem[1173] = 190;
razn_h_mem[1174] = 66;
razn_h_mem[1175] = 196;
razn_h_mem[1176] = 72;
razn_h_mem[1177] = 202;
razn_h_mem[1178] = 78;
razn_h_mem[1179] = 208;
razn_h_mem[1180] = 84;
razn_h_mem[1181] = 214;
razn_h_mem[1182] = 90;
razn_h_mem[1183] = 220;
razn_h_mem[1184] = 96;
razn_h_mem[1185] = 226;
razn_h_mem[1186] = 102;
razn_h_mem[1187] = 232;
razn_h_mem[1188] = 108;
razn_h_mem[1189] = 238;
razn_h_mem[1190] = 114;
razn_h_mem[1191] = 244;
razn_h_mem[1192] = 120;
razn_h_mem[1193] = 250;
razn_h_mem[1194] = 126;
razn_h_mem[1195] = 2;
razn_h_mem[1196] = 132;
razn_h_mem[1197] = 8;
razn_h_mem[1198] = 138;
razn_h_mem[1199] = 14;
razn_h_mem[1200] = 144;
razn_h_mem[1201] = 20;
razn_h_mem[1202] = 150;
razn_h_mem[1203] = 26;
razn_h_mem[1204] = 156;
razn_h_mem[1205] = 32;
razn_h_mem[1206] = 162;
razn_h_mem[1207] = 38;
razn_h_mem[1208] = 168;
razn_h_mem[1209] = 44;
razn_h_mem[1210] = 174;
razn_h_mem[1211] = 50;
razn_h_mem[1212] = 180;
razn_h_mem[1213] = 56;
razn_h_mem[1214] = 186;
razn_h_mem[1215] = 62;
razn_h_mem[1216] = 192;
razn_h_mem[1217] = 68;
razn_h_mem[1218] = 198;
razn_h_mem[1219] = 74;
razn_h_mem[1220] = 204;
razn_h_mem[1221] = 80;
razn_h_mem[1222] = 210;
razn_h_mem[1223] = 86;
razn_h_mem[1224] = 216;
razn_h_mem[1225] = 92;
razn_h_mem[1226] = 222;
razn_h_mem[1227] = 98;
razn_h_mem[1228] = 228;
razn_h_mem[1229] = 104;
razn_h_mem[1230] = 234;
razn_h_mem[1231] = 110;
razn_h_mem[1232] = 240;
razn_h_mem[1233] = 116;
razn_h_mem[1234] = 246;
razn_h_mem[1235] = 122;
razn_h_mem[1236] = 252;
razn_h_mem[1237] = 128;
razn_h_mem[1238] = 4;
razn_h_mem[1239] = 134;
razn_h_mem[1240] = 10;
razn_h_mem[1241] = 140;
razn_h_mem[1242] = 16;
razn_h_mem[1243] = 146;
razn_h_mem[1244] = 22;
razn_h_mem[1245] = 152;
razn_h_mem[1246] = 28;
razn_h_mem[1247] = 158;
razn_h_mem[1248] = 34;
razn_h_mem[1249] = 164;
razn_h_mem[1250] = 40;
razn_h_mem[1251] = 170;
razn_h_mem[1252] = 46;
razn_h_mem[1253] = 176;
razn_h_mem[1254] = 52;
razn_h_mem[1255] = 182;
razn_h_mem[1256] = 58;
razn_h_mem[1257] = 188;
razn_h_mem[1258] = 64;
razn_h_mem[1259] = 194;
razn_h_mem[1260] = 70;
razn_h_mem[1261] = 200;
razn_h_mem[1262] = 76;
razn_h_mem[1263] = 206;
razn_h_mem[1264] = 82;
razn_h_mem[1265] = 212;
razn_h_mem[1266] = 88;
razn_h_mem[1267] = 218;
razn_h_mem[1268] = 94;
razn_h_mem[1269] = 224;
razn_h_mem[1270] = 100;
razn_h_mem[1271] = 230;
razn_h_mem[1272] = 106;
razn_h_mem[1273] = 236;
razn_h_mem[1274] = 112;
razn_h_mem[1275] = 242;
razn_h_mem[1276] = 118;
razn_h_mem[1277] = 248;
razn_h_mem[1278] = 124;
razn_h_mem[1279] = 255;
razn_h_mem[1280] = 0;
razn_h_mem[1281] = 130;
razn_h_mem[1282] = 6;
razn_h_mem[1283] = 136;
razn_h_mem[1284] = 12;
razn_h_mem[1285] = 142;
razn_h_mem[1286] = 18;
razn_h_mem[1287] = 148;
razn_h_mem[1288] = 24;
razn_h_mem[1289] = 154;
razn_h_mem[1290] = 30;
razn_h_mem[1291] = 160;
razn_h_mem[1292] = 36;
razn_h_mem[1293] = 166;
razn_h_mem[1294] = 42;
razn_h_mem[1295] = 172;
razn_h_mem[1296] = 48;
razn_h_mem[1297] = 178;
razn_h_mem[1298] = 54;
razn_h_mem[1299] = 184;
razn_h_mem[1300] = 60;
razn_h_mem[1301] = 190;
razn_h_mem[1302] = 66;
razn_h_mem[1303] = 196;
razn_h_mem[1304] = 72;
razn_h_mem[1305] = 202;
razn_h_mem[1306] = 78;
razn_h_mem[1307] = 208;
razn_h_mem[1308] = 84;
razn_h_mem[1309] = 214;
razn_h_mem[1310] = 90;
razn_h_mem[1311] = 220;
razn_h_mem[1312] = 96;
razn_h_mem[1313] = 226;
razn_h_mem[1314] = 102;
razn_h_mem[1315] = 232;
razn_h_mem[1316] = 108;
razn_h_mem[1317] = 238;
razn_h_mem[1318] = 114;
razn_h_mem[1319] = 244;
razn_h_mem[1320] = 120;
razn_h_mem[1321] = 250;
razn_h_mem[1322] = 126;
razn_h_mem[1323] = 2;
razn_h_mem[1324] = 132;
razn_h_mem[1325] = 8;
razn_h_mem[1326] = 138;
razn_h_mem[1327] = 14;
razn_h_mem[1328] = 144;
razn_h_mem[1329] = 20;
razn_h_mem[1330] = 150;
razn_h_mem[1331] = 26;
razn_h_mem[1332] = 156;
razn_h_mem[1333] = 32;
razn_h_mem[1334] = 162;
razn_h_mem[1335] = 38;
razn_h_mem[1336] = 168;
razn_h_mem[1337] = 44;
razn_h_mem[1338] = 174;
razn_h_mem[1339] = 50;
razn_h_mem[1340] = 180;
razn_h_mem[1341] = 56;
razn_h_mem[1342] = 186;
razn_h_mem[1343] = 62;
razn_h_mem[1344] = 192;
razn_h_mem[1345] = 68;
razn_h_mem[1346] = 198;
razn_h_mem[1347] = 74;
razn_h_mem[1348] = 204;
razn_h_mem[1349] = 80;
razn_h_mem[1350] = 210;
razn_h_mem[1351] = 86;
razn_h_mem[1352] = 216;
razn_h_mem[1353] = 92;
razn_h_mem[1354] = 222;
razn_h_mem[1355] = 98;
razn_h_mem[1356] = 228;
razn_h_mem[1357] = 104;
razn_h_mem[1358] = 234;
razn_h_mem[1359] = 110;
razn_h_mem[1360] = 240;
razn_h_mem[1361] = 116;
razn_h_mem[1362] = 246;
razn_h_mem[1363] = 122;
razn_h_mem[1364] = 252;
razn_h_mem[1365] = 128;
razn_h_mem[1366] = 4;
razn_h_mem[1367] = 134;
razn_h_mem[1368] = 10;
razn_h_mem[1369] = 140;
razn_h_mem[1370] = 16;
razn_h_mem[1371] = 146;
razn_h_mem[1372] = 22;
razn_h_mem[1373] = 152;
razn_h_mem[1374] = 28;
razn_h_mem[1375] = 158;
razn_h_mem[1376] = 34;
razn_h_mem[1377] = 164;
razn_h_mem[1378] = 40;
razn_h_mem[1379] = 170;
razn_h_mem[1380] = 46;
razn_h_mem[1381] = 176;
razn_h_mem[1382] = 52;
razn_h_mem[1383] = 182;
razn_h_mem[1384] = 58;
razn_h_mem[1385] = 188;
razn_h_mem[1386] = 64;
razn_h_mem[1387] = 194;
razn_h_mem[1388] = 70;
razn_h_mem[1389] = 200;
razn_h_mem[1390] = 76;
razn_h_mem[1391] = 206;
razn_h_mem[1392] = 82;
razn_h_mem[1393] = 212;
razn_h_mem[1394] = 88;
razn_h_mem[1395] = 218;
razn_h_mem[1396] = 94;
razn_h_mem[1397] = 224;
razn_h_mem[1398] = 100;
razn_h_mem[1399] = 230;
razn_h_mem[1400] = 106;
razn_h_mem[1401] = 236;
razn_h_mem[1402] = 112;
razn_h_mem[1403] = 242;
razn_h_mem[1404] = 118;
razn_h_mem[1405] = 248;
razn_h_mem[1406] = 124;
razn_h_mem[1407] = 255;
razn_h_mem[1408] = 0;
razn_h_mem[1409] = 130;
razn_h_mem[1410] = 6;
razn_h_mem[1411] = 136;
razn_h_mem[1412] = 12;
razn_h_mem[1413] = 142;
razn_h_mem[1414] = 18;
razn_h_mem[1415] = 148;
razn_h_mem[1416] = 24;
razn_h_mem[1417] = 154;
razn_h_mem[1418] = 30;
razn_h_mem[1419] = 160;
razn_h_mem[1420] = 36;
razn_h_mem[1421] = 166;
razn_h_mem[1422] = 42;
razn_h_mem[1423] = 172;
razn_h_mem[1424] = 48;
razn_h_mem[1425] = 178;
razn_h_mem[1426] = 54;
razn_h_mem[1427] = 184;
razn_h_mem[1428] = 60;
razn_h_mem[1429] = 190;
razn_h_mem[1430] = 66;
razn_h_mem[1431] = 196;
razn_h_mem[1432] = 72;
razn_h_mem[1433] = 202;
razn_h_mem[1434] = 78;
razn_h_mem[1435] = 208;
razn_h_mem[1436] = 84;
razn_h_mem[1437] = 214;
razn_h_mem[1438] = 90;
razn_h_mem[1439] = 220;
razn_h_mem[1440] = 96;
razn_h_mem[1441] = 226;
razn_h_mem[1442] = 102;
razn_h_mem[1443] = 232;
razn_h_mem[1444] = 108;
razn_h_mem[1445] = 238;
razn_h_mem[1446] = 114;
razn_h_mem[1447] = 244;
razn_h_mem[1448] = 120;
razn_h_mem[1449] = 250;
razn_h_mem[1450] = 126;
razn_h_mem[1451] = 2;
razn_h_mem[1452] = 132;
razn_h_mem[1453] = 8;
razn_h_mem[1454] = 138;
razn_h_mem[1455] = 14;
razn_h_mem[1456] = 144;
razn_h_mem[1457] = 20;
razn_h_mem[1458] = 150;
razn_h_mem[1459] = 26;
razn_h_mem[1460] = 156;
razn_h_mem[1461] = 32;
razn_h_mem[1462] = 162;
razn_h_mem[1463] = 38;
razn_h_mem[1464] = 168;
razn_h_mem[1465] = 44;
razn_h_mem[1466] = 174;
razn_h_mem[1467] = 50;
razn_h_mem[1468] = 180;
razn_h_mem[1469] = 56;
razn_h_mem[1470] = 186;
razn_h_mem[1471] = 62;
razn_h_mem[1472] = 192;
razn_h_mem[1473] = 68;
razn_h_mem[1474] = 198;
razn_h_mem[1475] = 74;
razn_h_mem[1476] = 204;
razn_h_mem[1477] = 80;
razn_h_mem[1478] = 210;
razn_h_mem[1479] = 86;
razn_h_mem[1480] = 216;
razn_h_mem[1481] = 92;
razn_h_mem[1482] = 222;
razn_h_mem[1483] = 98;
razn_h_mem[1484] = 228;
razn_h_mem[1485] = 104;
razn_h_mem[1486] = 234;
razn_h_mem[1487] = 110;
razn_h_mem[1488] = 240;
razn_h_mem[1489] = 116;
razn_h_mem[1490] = 246;
razn_h_mem[1491] = 122;
razn_h_mem[1492] = 252;
razn_h_mem[1493] = 128;
razn_h_mem[1494] = 4;
razn_h_mem[1495] = 134;
razn_h_mem[1496] = 10;
razn_h_mem[1497] = 140;
razn_h_mem[1498] = 16;
razn_h_mem[1499] = 146;
razn_h_mem[1500] = 22;
razn_h_mem[1501] = 152;
razn_h_mem[1502] = 28;
razn_h_mem[1503] = 158;
razn_h_mem[1504] = 34;
razn_h_mem[1505] = 164;
razn_h_mem[1506] = 40;
razn_h_mem[1507] = 170;
razn_h_mem[1508] = 46;
razn_h_mem[1509] = 176;
razn_h_mem[1510] = 52;
razn_h_mem[1511] = 182;
razn_h_mem[1512] = 58;
razn_h_mem[1513] = 188;
razn_h_mem[1514] = 64;
razn_h_mem[1515] = 194;
razn_h_mem[1516] = 70;
razn_h_mem[1517] = 200;
razn_h_mem[1518] = 76;
razn_h_mem[1519] = 206;
razn_h_mem[1520] = 82;
razn_h_mem[1521] = 212;
razn_h_mem[1522] = 88;
razn_h_mem[1523] = 218;
razn_h_mem[1524] = 94;
razn_h_mem[1525] = 224;
razn_h_mem[1526] = 100;
razn_h_mem[1527] = 230;
razn_h_mem[1528] = 106;
razn_h_mem[1529] = 236;
razn_h_mem[1530] = 112;
razn_h_mem[1531] = 242;
razn_h_mem[1532] = 118;
razn_h_mem[1533] = 248;
razn_h_mem[1534] = 124;
razn_h_mem[1535] = 255;
razn_h_mem[1536] = 0;
razn_h_mem[1537] = 130;
razn_h_mem[1538] = 6;
razn_h_mem[1539] = 136;
razn_h_mem[1540] = 12;
razn_h_mem[1541] = 142;
razn_h_mem[1542] = 18;
razn_h_mem[1543] = 148;
razn_h_mem[1544] = 24;
razn_h_mem[1545] = 154;
razn_h_mem[1546] = 30;
razn_h_mem[1547] = 160;
razn_h_mem[1548] = 36;
razn_h_mem[1549] = 166;
razn_h_mem[1550] = 42;
razn_h_mem[1551] = 172;
razn_h_mem[1552] = 48;
razn_h_mem[1553] = 178;
razn_h_mem[1554] = 54;
razn_h_mem[1555] = 184;
razn_h_mem[1556] = 60;
razn_h_mem[1557] = 190;
razn_h_mem[1558] = 66;
razn_h_mem[1559] = 196;
razn_h_mem[1560] = 72;
razn_h_mem[1561] = 202;
razn_h_mem[1562] = 78;
razn_h_mem[1563] = 208;
razn_h_mem[1564] = 84;
razn_h_mem[1565] = 214;
razn_h_mem[1566] = 90;
razn_h_mem[1567] = 220;
razn_h_mem[1568] = 96;
razn_h_mem[1569] = 226;
razn_h_mem[1570] = 102;
razn_h_mem[1571] = 232;
razn_h_mem[1572] = 108;
razn_h_mem[1573] = 238;
razn_h_mem[1574] = 114;
razn_h_mem[1575] = 244;
razn_h_mem[1576] = 120;
razn_h_mem[1577] = 250;
razn_h_mem[1578] = 126;
razn_h_mem[1579] = 2;
razn_h_mem[1580] = 132;
razn_h_mem[1581] = 8;
razn_h_mem[1582] = 138;
razn_h_mem[1583] = 14;
razn_h_mem[1584] = 144;
razn_h_mem[1585] = 20;
razn_h_mem[1586] = 150;
razn_h_mem[1587] = 26;
razn_h_mem[1588] = 156;
razn_h_mem[1589] = 32;
razn_h_mem[1590] = 162;
razn_h_mem[1591] = 38;
razn_h_mem[1592] = 168;
razn_h_mem[1593] = 44;
razn_h_mem[1594] = 174;
razn_h_mem[1595] = 50;
razn_h_mem[1596] = 180;
razn_h_mem[1597] = 56;
razn_h_mem[1598] = 186;
razn_h_mem[1599] = 62;
razn_h_mem[1600] = 192;
razn_h_mem[1601] = 68;
razn_h_mem[1602] = 198;
razn_h_mem[1603] = 74;
razn_h_mem[1604] = 204;
razn_h_mem[1605] = 80;
razn_h_mem[1606] = 210;
razn_h_mem[1607] = 86;
razn_h_mem[1608] = 216;
razn_h_mem[1609] = 92;
razn_h_mem[1610] = 222;
razn_h_mem[1611] = 98;
razn_h_mem[1612] = 228;
razn_h_mem[1613] = 104;
razn_h_mem[1614] = 234;
razn_h_mem[1615] = 110;
razn_h_mem[1616] = 240;
razn_h_mem[1617] = 116;
razn_h_mem[1618] = 246;
razn_h_mem[1619] = 122;
razn_h_mem[1620] = 252;
razn_h_mem[1621] = 128;
razn_h_mem[1622] = 4;
razn_h_mem[1623] = 134;
razn_h_mem[1624] = 10;
razn_h_mem[1625] = 140;
razn_h_mem[1626] = 16;
razn_h_mem[1627] = 146;
razn_h_mem[1628] = 22;
razn_h_mem[1629] = 152;
razn_h_mem[1630] = 28;
razn_h_mem[1631] = 158;
razn_h_mem[1632] = 34;
razn_h_mem[1633] = 164;
razn_h_mem[1634] = 40;
razn_h_mem[1635] = 170;
razn_h_mem[1636] = 46;
razn_h_mem[1637] = 176;
razn_h_mem[1638] = 52;
razn_h_mem[1639] = 182;
razn_h_mem[1640] = 58;
razn_h_mem[1641] = 188;
razn_h_mem[1642] = 64;
razn_h_mem[1643] = 194;
razn_h_mem[1644] = 70;
razn_h_mem[1645] = 200;
razn_h_mem[1646] = 76;
razn_h_mem[1647] = 206;
razn_h_mem[1648] = 82;
razn_h_mem[1649] = 212;
razn_h_mem[1650] = 88;
razn_h_mem[1651] = 218;
razn_h_mem[1652] = 94;
razn_h_mem[1653] = 224;
razn_h_mem[1654] = 100;
razn_h_mem[1655] = 230;
razn_h_mem[1656] = 106;
razn_h_mem[1657] = 236;
razn_h_mem[1658] = 112;
razn_h_mem[1659] = 242;
razn_h_mem[1660] = 118;
razn_h_mem[1661] = 248;
razn_h_mem[1662] = 124;
razn_h_mem[1663] = 255;
razn_h_mem[1664] = 0;
razn_h_mem[1665] = 130;
razn_h_mem[1666] = 6;
razn_h_mem[1667] = 136;
razn_h_mem[1668] = 12;
razn_h_mem[1669] = 142;
razn_h_mem[1670] = 18;
razn_h_mem[1671] = 148;
razn_h_mem[1672] = 24;
razn_h_mem[1673] = 154;
razn_h_mem[1674] = 30;
razn_h_mem[1675] = 160;
razn_h_mem[1676] = 36;
razn_h_mem[1677] = 166;
razn_h_mem[1678] = 42;
razn_h_mem[1679] = 172;
razn_h_mem[1680] = 48;
razn_h_mem[1681] = 178;
razn_h_mem[1682] = 54;
razn_h_mem[1683] = 184;
razn_h_mem[1684] = 60;
razn_h_mem[1685] = 190;
razn_h_mem[1686] = 66;
razn_h_mem[1687] = 196;
razn_h_mem[1688] = 72;
razn_h_mem[1689] = 202;
razn_h_mem[1690] = 78;
razn_h_mem[1691] = 208;
razn_h_mem[1692] = 84;
razn_h_mem[1693] = 214;
razn_h_mem[1694] = 90;
razn_h_mem[1695] = 220;
razn_h_mem[1696] = 96;
razn_h_mem[1697] = 226;
razn_h_mem[1698] = 102;
razn_h_mem[1699] = 232;
razn_h_mem[1700] = 108;
razn_h_mem[1701] = 238;
razn_h_mem[1702] = 114;
razn_h_mem[1703] = 244;
razn_h_mem[1704] = 120;
razn_h_mem[1705] = 250;
razn_h_mem[1706] = 126;
razn_h_mem[1707] = 2;
razn_h_mem[1708] = 132;
razn_h_mem[1709] = 8;
razn_h_mem[1710] = 138;
razn_h_mem[1711] = 14;
razn_h_mem[1712] = 144;
razn_h_mem[1713] = 20;
razn_h_mem[1714] = 150;
razn_h_mem[1715] = 26;
razn_h_mem[1716] = 156;
razn_h_mem[1717] = 32;
razn_h_mem[1718] = 162;
razn_h_mem[1719] = 38;
razn_h_mem[1720] = 168;
razn_h_mem[1721] = 44;
razn_h_mem[1722] = 174;
razn_h_mem[1723] = 50;
razn_h_mem[1724] = 180;
razn_h_mem[1725] = 56;
razn_h_mem[1726] = 186;
razn_h_mem[1727] = 62;
razn_h_mem[1728] = 192;
razn_h_mem[1729] = 68;
razn_h_mem[1730] = 198;
razn_h_mem[1731] = 74;
razn_h_mem[1732] = 204;
razn_h_mem[1733] = 80;
razn_h_mem[1734] = 210;
razn_h_mem[1735] = 86;
razn_h_mem[1736] = 216;
razn_h_mem[1737] = 92;
razn_h_mem[1738] = 222;
razn_h_mem[1739] = 98;
razn_h_mem[1740] = 228;
razn_h_mem[1741] = 104;
razn_h_mem[1742] = 234;
razn_h_mem[1743] = 110;
razn_h_mem[1744] = 240;
razn_h_mem[1745] = 116;
razn_h_mem[1746] = 246;
razn_h_mem[1747] = 122;
razn_h_mem[1748] = 252;
razn_h_mem[1749] = 128;
razn_h_mem[1750] = 4;
razn_h_mem[1751] = 134;
razn_h_mem[1752] = 10;
razn_h_mem[1753] = 140;
razn_h_mem[1754] = 16;
razn_h_mem[1755] = 146;
razn_h_mem[1756] = 22;
razn_h_mem[1757] = 152;
razn_h_mem[1758] = 28;
razn_h_mem[1759] = 158;
razn_h_mem[1760] = 34;
razn_h_mem[1761] = 164;
razn_h_mem[1762] = 40;
razn_h_mem[1763] = 170;
razn_h_mem[1764] = 46;
razn_h_mem[1765] = 176;
razn_h_mem[1766] = 52;
razn_h_mem[1767] = 182;
razn_h_mem[1768] = 58;
razn_h_mem[1769] = 188;
razn_h_mem[1770] = 64;
razn_h_mem[1771] = 194;
razn_h_mem[1772] = 70;
razn_h_mem[1773] = 200;
razn_h_mem[1774] = 76;
razn_h_mem[1775] = 206;
razn_h_mem[1776] = 82;
razn_h_mem[1777] = 212;
razn_h_mem[1778] = 88;
razn_h_mem[1779] = 218;
razn_h_mem[1780] = 94;
razn_h_mem[1781] = 224;
razn_h_mem[1782] = 100;
razn_h_mem[1783] = 230;
razn_h_mem[1784] = 106;
razn_h_mem[1785] = 236;
razn_h_mem[1786] = 112;
razn_h_mem[1787] = 242;
razn_h_mem[1788] = 118;
razn_h_mem[1789] = 248;
razn_h_mem[1790] = 124;
razn_h_mem[1791] = 255;
razn_h_mem[1792] = 0;
razn_h_mem[1793] = 130;
razn_h_mem[1794] = 6;
razn_h_mem[1795] = 136;
razn_h_mem[1796] = 12;
razn_h_mem[1797] = 142;
razn_h_mem[1798] = 18;
razn_h_mem[1799] = 148;
razn_h_mem[1800] = 24;
razn_h_mem[1801] = 154;
razn_h_mem[1802] = 30;
razn_h_mem[1803] = 160;
razn_h_mem[1804] = 36;
razn_h_mem[1805] = 166;
razn_h_mem[1806] = 42;
razn_h_mem[1807] = 172;
razn_h_mem[1808] = 48;
razn_h_mem[1809] = 178;
razn_h_mem[1810] = 54;
razn_h_mem[1811] = 184;
razn_h_mem[1812] = 60;
razn_h_mem[1813] = 190;
razn_h_mem[1814] = 66;
razn_h_mem[1815] = 196;
razn_h_mem[1816] = 72;
razn_h_mem[1817] = 202;
razn_h_mem[1818] = 78;
razn_h_mem[1819] = 208;
razn_h_mem[1820] = 84;
razn_h_mem[1821] = 214;
razn_h_mem[1822] = 90;
razn_h_mem[1823] = 220;
razn_h_mem[1824] = 96;
razn_h_mem[1825] = 226;
razn_h_mem[1826] = 102;
razn_h_mem[1827] = 232;
razn_h_mem[1828] = 108;
razn_h_mem[1829] = 238;
razn_h_mem[1830] = 114;
razn_h_mem[1831] = 244;
razn_h_mem[1832] = 120;
razn_h_mem[1833] = 250;
razn_h_mem[1834] = 126;
razn_h_mem[1835] = 2;
razn_h_mem[1836] = 132;
razn_h_mem[1837] = 8;
razn_h_mem[1838] = 138;
razn_h_mem[1839] = 14;
razn_h_mem[1840] = 144;
razn_h_mem[1841] = 20;
razn_h_mem[1842] = 150;
razn_h_mem[1843] = 26;
razn_h_mem[1844] = 156;
razn_h_mem[1845] = 32;
razn_h_mem[1846] = 162;
razn_h_mem[1847] = 38;
razn_h_mem[1848] = 168;
razn_h_mem[1849] = 44;
razn_h_mem[1850] = 174;
razn_h_mem[1851] = 50;
razn_h_mem[1852] = 180;
razn_h_mem[1853] = 56;
razn_h_mem[1854] = 186;
razn_h_mem[1855] = 62;
razn_h_mem[1856] = 192;
razn_h_mem[1857] = 68;
razn_h_mem[1858] = 198;
razn_h_mem[1859] = 74;
razn_h_mem[1860] = 204;
razn_h_mem[1861] = 80;
razn_h_mem[1862] = 210;
razn_h_mem[1863] = 86;
razn_h_mem[1864] = 216;
razn_h_mem[1865] = 92;
razn_h_mem[1866] = 222;
razn_h_mem[1867] = 98;
razn_h_mem[1868] = 228;
razn_h_mem[1869] = 104;
razn_h_mem[1870] = 234;
razn_h_mem[1871] = 110;
razn_h_mem[1872] = 240;
razn_h_mem[1873] = 116;
razn_h_mem[1874] = 246;
razn_h_mem[1875] = 122;
razn_h_mem[1876] = 252;
razn_h_mem[1877] = 128;
razn_h_mem[1878] = 4;
razn_h_mem[1879] = 134;
razn_h_mem[1880] = 10;
razn_h_mem[1881] = 140;
razn_h_mem[1882] = 16;
razn_h_mem[1883] = 146;
razn_h_mem[1884] = 22;
razn_h_mem[1885] = 152;
razn_h_mem[1886] = 28;
razn_h_mem[1887] = 158;
razn_h_mem[1888] = 34;
razn_h_mem[1889] = 164;
razn_h_mem[1890] = 40;
razn_h_mem[1891] = 170;
razn_h_mem[1892] = 46;
razn_h_mem[1893] = 176;
razn_h_mem[1894] = 52;
razn_h_mem[1895] = 182;
razn_h_mem[1896] = 58;
razn_h_mem[1897] = 188;
razn_h_mem[1898] = 64;
razn_h_mem[1899] = 194;
razn_h_mem[1900] = 70;
razn_h_mem[1901] = 200;
razn_h_mem[1902] = 76;
razn_h_mem[1903] = 206;
razn_h_mem[1904] = 82;
razn_h_mem[1905] = 212;
razn_h_mem[1906] = 88;
razn_h_mem[1907] = 218;
razn_h_mem[1908] = 94;
razn_h_mem[1909] = 224;
razn_h_mem[1910] = 100;
razn_h_mem[1911] = 230;
razn_h_mem[1912] = 106;
razn_h_mem[1913] = 236;
razn_h_mem[1914] = 112;
razn_h_mem[1915] = 242;
razn_h_mem[1916] = 118;
razn_h_mem[1917] = 248;
razn_h_mem[1918] = 124;
razn_h_mem[1919] = 255;
razn_h_mem[1920] = 0;
razn_h_mem[1921] = 130;
razn_h_mem[1922] = 6;
razn_h_mem[1923] = 136;
razn_h_mem[1924] = 12;
razn_h_mem[1925] = 142;
razn_h_mem[1926] = 18;
razn_h_mem[1927] = 148;
razn_h_mem[1928] = 24;
razn_h_mem[1929] = 154;
razn_h_mem[1930] = 30;
razn_h_mem[1931] = 160;
razn_h_mem[1932] = 36;
razn_h_mem[1933] = 166;
razn_h_mem[1934] = 42;
razn_h_mem[1935] = 172;
razn_h_mem[1936] = 48;
razn_h_mem[1937] = 178;
razn_h_mem[1938] = 54;
razn_h_mem[1939] = 184;
razn_h_mem[1940] = 60;
razn_h_mem[1941] = 190;
razn_h_mem[1942] = 66;
razn_h_mem[1943] = 196;
razn_h_mem[1944] = 72;
razn_h_mem[1945] = 202;
razn_h_mem[1946] = 78;
razn_h_mem[1947] = 208;
razn_h_mem[1948] = 84;
razn_h_mem[1949] = 214;
razn_h_mem[1950] = 90;
razn_h_mem[1951] = 220;
razn_h_mem[1952] = 96;
razn_h_mem[1953] = 226;
razn_h_mem[1954] = 102;
razn_h_mem[1955] = 232;
razn_h_mem[1956] = 108;
razn_h_mem[1957] = 238;
razn_h_mem[1958] = 114;
razn_h_mem[1959] = 244;
razn_h_mem[1960] = 120;
razn_h_mem[1961] = 250;
razn_h_mem[1962] = 126;
razn_h_mem[1963] = 2;
razn_h_mem[1964] = 132;
razn_h_mem[1965] = 8;
razn_h_mem[1966] = 138;
razn_h_mem[1967] = 14;
razn_h_mem[1968] = 144;
razn_h_mem[1969] = 20;
razn_h_mem[1970] = 150;
razn_h_mem[1971] = 26;
razn_h_mem[1972] = 156;
razn_h_mem[1973] = 32;
razn_h_mem[1974] = 162;
razn_h_mem[1975] = 38;
razn_h_mem[1976] = 168;
razn_h_mem[1977] = 44;
razn_h_mem[1978] = 174;
razn_h_mem[1979] = 50;
razn_h_mem[1980] = 180;
razn_h_mem[1981] = 56;
razn_h_mem[1982] = 186;
razn_h_mem[1983] = 62;
razn_h_mem[1984] = 192;
razn_h_mem[1985] = 68;
razn_h_mem[1986] = 198;
razn_h_mem[1987] = 74;
razn_h_mem[1988] = 204;
razn_h_mem[1989] = 80;
razn_h_mem[1990] = 210;
razn_h_mem[1991] = 86;
razn_h_mem[1992] = 216;
razn_h_mem[1993] = 92;
razn_h_mem[1994] = 222;
razn_h_mem[1995] = 98;
razn_h_mem[1996] = 228;
razn_h_mem[1997] = 104;
razn_h_mem[1998] = 234;
razn_h_mem[1999] = 110;
razn_h_mem[2000] = 240;
razn_h_mem[2001] = 116;
razn_h_mem[2002] = 246;
razn_h_mem[2003] = 122;
razn_h_mem[2004] = 252;
razn_h_mem[2005] = 128;
razn_h_mem[2006] = 4;
razn_h_mem[2007] = 134;
razn_h_mem[2008] = 10;
razn_h_mem[2009] = 140;
razn_h_mem[2010] = 16;
razn_h_mem[2011] = 146;
razn_h_mem[2012] = 22;
razn_h_mem[2013] = 152;
razn_h_mem[2014] = 28;
razn_h_mem[2015] = 158;
razn_h_mem[2016] = 34;
razn_h_mem[2017] = 164;
razn_h_mem[2018] = 40;
razn_h_mem[2019] = 170;
razn_h_mem[2020] = 46;
razn_h_mem[2021] = 176;
razn_h_mem[2022] = 52;
razn_h_mem[2023] = 182;
razn_h_mem[2024] = 58;
razn_h_mem[2025] = 188;
razn_h_mem[2026] = 64;
razn_h_mem[2027] = 194;
razn_h_mem[2028] = 70;
razn_h_mem[2029] = 200;
razn_h_mem[2030] = 76;
razn_h_mem[2031] = 206;
razn_h_mem[2032] = 82;
razn_h_mem[2033] = 212;
razn_h_mem[2034] = 88;
razn_h_mem[2035] = 218;
razn_h_mem[2036] = 94;
razn_h_mem[2037] = 224;
razn_h_mem[2038] = 100;
razn_h_mem[2039] = 230;
razn_h_mem[2040] = 106;
razn_h_mem[2041] = 236;
razn_h_mem[2042] = 112;
razn_h_mem[2043] = 242;
razn_h_mem[2044] = 118;
razn_h_mem[2045] = 248;
razn_h_mem[2046] = 124;
razn_h_mem[2047] = 255;
razn_h_mem[2048] = 0;
razn_h_mem[2049] = 130;
razn_h_mem[2050] = 6;
razn_h_mem[2051] = 136;
razn_h_mem[2052] = 12;
razn_h_mem[2053] = 142;
razn_h_mem[2054] = 18;
razn_h_mem[2055] = 148;
razn_h_mem[2056] = 24;
razn_h_mem[2057] = 154;
razn_h_mem[2058] = 30;
razn_h_mem[2059] = 160;
razn_h_mem[2060] = 36;
razn_h_mem[2061] = 166;
razn_h_mem[2062] = 42;
razn_h_mem[2063] = 172;
razn_h_mem[2064] = 48;
razn_h_mem[2065] = 178;
razn_h_mem[2066] = 54;
razn_h_mem[2067] = 184;
razn_h_mem[2068] = 60;
razn_h_mem[2069] = 190;
razn_h_mem[2070] = 66;
razn_h_mem[2071] = 196;
razn_h_mem[2072] = 72;
razn_h_mem[2073] = 202;
razn_h_mem[2074] = 78;
razn_h_mem[2075] = 208;
razn_h_mem[2076] = 84;
razn_h_mem[2077] = 214;
razn_h_mem[2078] = 90;
razn_h_mem[2079] = 220;
razn_h_mem[2080] = 96;
razn_h_mem[2081] = 226;
razn_h_mem[2082] = 102;
razn_h_mem[2083] = 232;
razn_h_mem[2084] = 108;
razn_h_mem[2085] = 238;
razn_h_mem[2086] = 114;
razn_h_mem[2087] = 244;
razn_h_mem[2088] = 120;
razn_h_mem[2089] = 250;
razn_h_mem[2090] = 126;
razn_h_mem[2091] = 2;
razn_h_mem[2092] = 132;
razn_h_mem[2093] = 8;
razn_h_mem[2094] = 138;
razn_h_mem[2095] = 14;
razn_h_mem[2096] = 144;
razn_h_mem[2097] = 20;
razn_h_mem[2098] = 150;
razn_h_mem[2099] = 26;
razn_h_mem[2100] = 156;
razn_h_mem[2101] = 32;
razn_h_mem[2102] = 162;
razn_h_mem[2103] = 38;
razn_h_mem[2104] = 168;
razn_h_mem[2105] = 44;
razn_h_mem[2106] = 174;
razn_h_mem[2107] = 50;
razn_h_mem[2108] = 180;
razn_h_mem[2109] = 56;
razn_h_mem[2110] = 186;
razn_h_mem[2111] = 62;
razn_h_mem[2112] = 192;
razn_h_mem[2113] = 68;
razn_h_mem[2114] = 198;
razn_h_mem[2115] = 74;
razn_h_mem[2116] = 204;
razn_h_mem[2117] = 80;
razn_h_mem[2118] = 210;
razn_h_mem[2119] = 86;
razn_h_mem[2120] = 216;
razn_h_mem[2121] = 92;
razn_h_mem[2122] = 222;
razn_h_mem[2123] = 98;
razn_h_mem[2124] = 228;
razn_h_mem[2125] = 104;
razn_h_mem[2126] = 234;
razn_h_mem[2127] = 110;
razn_h_mem[2128] = 240;
razn_h_mem[2129] = 116;
razn_h_mem[2130] = 246;
razn_h_mem[2131] = 122;
razn_h_mem[2132] = 252;
razn_h_mem[2133] = 128;
razn_h_mem[2134] = 4;
razn_h_mem[2135] = 134;
razn_h_mem[2136] = 10;
razn_h_mem[2137] = 140;
razn_h_mem[2138] = 16;
razn_h_mem[2139] = 146;
razn_h_mem[2140] = 22;
razn_h_mem[2141] = 152;
razn_h_mem[2142] = 28;
razn_h_mem[2143] = 158;
razn_h_mem[2144] = 34;
razn_h_mem[2145] = 164;
razn_h_mem[2146] = 40;
razn_h_mem[2147] = 170;
razn_h_mem[2148] = 46;
razn_h_mem[2149] = 176;
razn_h_mem[2150] = 52;
razn_h_mem[2151] = 182;
razn_h_mem[2152] = 58;
razn_h_mem[2153] = 188;
razn_h_mem[2154] = 64;
razn_h_mem[2155] = 194;
razn_h_mem[2156] = 70;
razn_h_mem[2157] = 200;
razn_h_mem[2158] = 76;
razn_h_mem[2159] = 206;
razn_h_mem[2160] = 82;
razn_h_mem[2161] = 212;
razn_h_mem[2162] = 88;
razn_h_mem[2163] = 218;
razn_h_mem[2164] = 94;
razn_h_mem[2165] = 224;
razn_h_mem[2166] = 100;
razn_h_mem[2167] = 230;
razn_h_mem[2168] = 106;
razn_h_mem[2169] = 236;
razn_h_mem[2170] = 112;
razn_h_mem[2171] = 242;
razn_h_mem[2172] = 118;
razn_h_mem[2173] = 248;
razn_h_mem[2174] = 124;
razn_h_mem[2175] = 255;
razn_h_mem[2176] = 0;
razn_h_mem[2177] = 130;
razn_h_mem[2178] = 6;
razn_h_mem[2179] = 136;
razn_h_mem[2180] = 12;
razn_h_mem[2181] = 142;
razn_h_mem[2182] = 18;
razn_h_mem[2183] = 148;
razn_h_mem[2184] = 24;
razn_h_mem[2185] = 154;
razn_h_mem[2186] = 30;
razn_h_mem[2187] = 160;
razn_h_mem[2188] = 36;
razn_h_mem[2189] = 166;
razn_h_mem[2190] = 42;
razn_h_mem[2191] = 172;
razn_h_mem[2192] = 48;
razn_h_mem[2193] = 178;
razn_h_mem[2194] = 54;
razn_h_mem[2195] = 184;
razn_h_mem[2196] = 60;
razn_h_mem[2197] = 190;
razn_h_mem[2198] = 66;
razn_h_mem[2199] = 196;
razn_h_mem[2200] = 72;
razn_h_mem[2201] = 202;
razn_h_mem[2202] = 78;
razn_h_mem[2203] = 208;
razn_h_mem[2204] = 84;
razn_h_mem[2205] = 214;
razn_h_mem[2206] = 90;
razn_h_mem[2207] = 220;
razn_h_mem[2208] = 96;
razn_h_mem[2209] = 226;
razn_h_mem[2210] = 102;
razn_h_mem[2211] = 232;
razn_h_mem[2212] = 108;
razn_h_mem[2213] = 238;
razn_h_mem[2214] = 114;
razn_h_mem[2215] = 244;
razn_h_mem[2216] = 120;
razn_h_mem[2217] = 250;
razn_h_mem[2218] = 126;
razn_h_mem[2219] = 2;
razn_h_mem[2220] = 132;
razn_h_mem[2221] = 8;
razn_h_mem[2222] = 138;
razn_h_mem[2223] = 14;
razn_h_mem[2224] = 144;
razn_h_mem[2225] = 20;
razn_h_mem[2226] = 150;
razn_h_mem[2227] = 26;
razn_h_mem[2228] = 156;
razn_h_mem[2229] = 32;
razn_h_mem[2230] = 162;
razn_h_mem[2231] = 38;
razn_h_mem[2232] = 168;
razn_h_mem[2233] = 44;
razn_h_mem[2234] = 174;
razn_h_mem[2235] = 50;
razn_h_mem[2236] = 180;
razn_h_mem[2237] = 56;
razn_h_mem[2238] = 186;
razn_h_mem[2239] = 62;
razn_h_mem[2240] = 192;
razn_h_mem[2241] = 68;
razn_h_mem[2242] = 198;
razn_h_mem[2243] = 74;
razn_h_mem[2244] = 204;
razn_h_mem[2245] = 80;
razn_h_mem[2246] = 210;
razn_h_mem[2247] = 86;
razn_h_mem[2248] = 216;
razn_h_mem[2249] = 92;
razn_h_mem[2250] = 222;
razn_h_mem[2251] = 98;
razn_h_mem[2252] = 228;
razn_h_mem[2253] = 104;
razn_h_mem[2254] = 234;
razn_h_mem[2255] = 110;
razn_h_mem[2256] = 240;
razn_h_mem[2257] = 116;
razn_h_mem[2258] = 246;
razn_h_mem[2259] = 122;
razn_h_mem[2260] = 252;
razn_h_mem[2261] = 128;
razn_h_mem[2262] = 4;
razn_h_mem[2263] = 134;
razn_h_mem[2264] = 10;
razn_h_mem[2265] = 140;
razn_h_mem[2266] = 16;
razn_h_mem[2267] = 146;
razn_h_mem[2268] = 22;
razn_h_mem[2269] = 152;
razn_h_mem[2270] = 28;
razn_h_mem[2271] = 158;
razn_h_mem[2272] = 34;
razn_h_mem[2273] = 164;
razn_h_mem[2274] = 40;
razn_h_mem[2275] = 170;
razn_h_mem[2276] = 46;
razn_h_mem[2277] = 176;
razn_h_mem[2278] = 52;
razn_h_mem[2279] = 182;
razn_h_mem[2280] = 58;
razn_h_mem[2281] = 188;
razn_h_mem[2282] = 64;
razn_h_mem[2283] = 194;
razn_h_mem[2284] = 70;
razn_h_mem[2285] = 200;
razn_h_mem[2286] = 76;
razn_h_mem[2287] = 206;
razn_h_mem[2288] = 82;
razn_h_mem[2289] = 212;
razn_h_mem[2290] = 88;
razn_h_mem[2291] = 218;
razn_h_mem[2292] = 94;
razn_h_mem[2293] = 224;
razn_h_mem[2294] = 100;
razn_h_mem[2295] = 230;
razn_h_mem[2296] = 106;
razn_h_mem[2297] = 236;
razn_h_mem[2298] = 112;
razn_h_mem[2299] = 242;
razn_h_mem[2300] = 118;
razn_h_mem[2301] = 248;
razn_h_mem[2302] = 124;
razn_h_mem[2303] = 255;
razn_h_mem[2304] = 0;
razn_h_mem[2305] = 130;
razn_h_mem[2306] = 6;
razn_h_mem[2307] = 136;
razn_h_mem[2308] = 12;
razn_h_mem[2309] = 142;
razn_h_mem[2310] = 18;
razn_h_mem[2311] = 148;
razn_h_mem[2312] = 24;
razn_h_mem[2313] = 154;
razn_h_mem[2314] = 30;
razn_h_mem[2315] = 160;
razn_h_mem[2316] = 36;
razn_h_mem[2317] = 166;
razn_h_mem[2318] = 42;
razn_h_mem[2319] = 172;
razn_h_mem[2320] = 48;
razn_h_mem[2321] = 178;
razn_h_mem[2322] = 54;
razn_h_mem[2323] = 184;
razn_h_mem[2324] = 60;
razn_h_mem[2325] = 190;
razn_h_mem[2326] = 66;
razn_h_mem[2327] = 196;
razn_h_mem[2328] = 72;
razn_h_mem[2329] = 202;
razn_h_mem[2330] = 78;
razn_h_mem[2331] = 208;
razn_h_mem[2332] = 84;
razn_h_mem[2333] = 214;
razn_h_mem[2334] = 90;
razn_h_mem[2335] = 220;
razn_h_mem[2336] = 96;
razn_h_mem[2337] = 226;
razn_h_mem[2338] = 102;
razn_h_mem[2339] = 232;
razn_h_mem[2340] = 108;
razn_h_mem[2341] = 238;
razn_h_mem[2342] = 114;
razn_h_mem[2343] = 244;
razn_h_mem[2344] = 120;
razn_h_mem[2345] = 250;
razn_h_mem[2346] = 126;
razn_h_mem[2347] = 2;
razn_h_mem[2348] = 132;
razn_h_mem[2349] = 8;
razn_h_mem[2350] = 138;
razn_h_mem[2351] = 14;
razn_h_mem[2352] = 144;
razn_h_mem[2353] = 20;
razn_h_mem[2354] = 150;
razn_h_mem[2355] = 26;
razn_h_mem[2356] = 156;
razn_h_mem[2357] = 32;
razn_h_mem[2358] = 162;
razn_h_mem[2359] = 38;
razn_h_mem[2360] = 168;
razn_h_mem[2361] = 44;
razn_h_mem[2362] = 174;
razn_h_mem[2363] = 50;
razn_h_mem[2364] = 180;
razn_h_mem[2365] = 56;
razn_h_mem[2366] = 186;
razn_h_mem[2367] = 62;
razn_h_mem[2368] = 192;
razn_h_mem[2369] = 68;
razn_h_mem[2370] = 198;
razn_h_mem[2371] = 74;
razn_h_mem[2372] = 204;
razn_h_mem[2373] = 80;
razn_h_mem[2374] = 210;
razn_h_mem[2375] = 86;
razn_h_mem[2376] = 216;
razn_h_mem[2377] = 92;
razn_h_mem[2378] = 222;
razn_h_mem[2379] = 98;
razn_h_mem[2380] = 228;
razn_h_mem[2381] = 104;
razn_h_mem[2382] = 234;
razn_h_mem[2383] = 110;
razn_h_mem[2384] = 240;
razn_h_mem[2385] = 116;
razn_h_mem[2386] = 246;
razn_h_mem[2387] = 122;
razn_h_mem[2388] = 252;
razn_h_mem[2389] = 128;
razn_h_mem[2390] = 4;
razn_h_mem[2391] = 134;
razn_h_mem[2392] = 10;
razn_h_mem[2393] = 140;
razn_h_mem[2394] = 16;
razn_h_mem[2395] = 146;
razn_h_mem[2396] = 22;
razn_h_mem[2397] = 152;
razn_h_mem[2398] = 28;
razn_h_mem[2399] = 158;
razn_h_mem[2400] = 34;
razn_h_mem[2401] = 164;
razn_h_mem[2402] = 40;
razn_h_mem[2403] = 170;
razn_h_mem[2404] = 46;
razn_h_mem[2405] = 176;
razn_h_mem[2406] = 52;
razn_h_mem[2407] = 182;
razn_h_mem[2408] = 58;
razn_h_mem[2409] = 188;
razn_h_mem[2410] = 64;
razn_h_mem[2411] = 194;
razn_h_mem[2412] = 70;
razn_h_mem[2413] = 200;
razn_h_mem[2414] = 76;
razn_h_mem[2415] = 206;
razn_h_mem[2416] = 82;
razn_h_mem[2417] = 212;
razn_h_mem[2418] = 88;
razn_h_mem[2419] = 218;
razn_h_mem[2420] = 94;
razn_h_mem[2421] = 224;
razn_h_mem[2422] = 100;
razn_h_mem[2423] = 230;
razn_h_mem[2424] = 106;
razn_h_mem[2425] = 236;
razn_h_mem[2426] = 112;
razn_h_mem[2427] = 242;
razn_h_mem[2428] = 118;
razn_h_mem[2429] = 248;
razn_h_mem[2430] = 124;
razn_h_mem[2431] = 255;
razn_h_mem[2432] = 0;
razn_h_mem[2433] = 130;
razn_h_mem[2434] = 6;
razn_h_mem[2435] = 136;
razn_h_mem[2436] = 12;
razn_h_mem[2437] = 142;
razn_h_mem[2438] = 18;
razn_h_mem[2439] = 148;
razn_h_mem[2440] = 24;
razn_h_mem[2441] = 154;
razn_h_mem[2442] = 30;
razn_h_mem[2443] = 160;
razn_h_mem[2444] = 36;
razn_h_mem[2445] = 166;
razn_h_mem[2446] = 42;
razn_h_mem[2447] = 172;
razn_h_mem[2448] = 48;
razn_h_mem[2449] = 178;
razn_h_mem[2450] = 54;
razn_h_mem[2451] = 184;
razn_h_mem[2452] = 60;
razn_h_mem[2453] = 190;
razn_h_mem[2454] = 66;
razn_h_mem[2455] = 196;
razn_h_mem[2456] = 72;
razn_h_mem[2457] = 202;
razn_h_mem[2458] = 78;
razn_h_mem[2459] = 208;
razn_h_mem[2460] = 84;
razn_h_mem[2461] = 214;
razn_h_mem[2462] = 90;
razn_h_mem[2463] = 220;
razn_h_mem[2464] = 96;
razn_h_mem[2465] = 226;
razn_h_mem[2466] = 102;
razn_h_mem[2467] = 232;
razn_h_mem[2468] = 108;
razn_h_mem[2469] = 238;
razn_h_mem[2470] = 114;
razn_h_mem[2471] = 244;
razn_h_mem[2472] = 120;
razn_h_mem[2473] = 250;
razn_h_mem[2474] = 126;
razn_h_mem[2475] = 2;
razn_h_mem[2476] = 132;
razn_h_mem[2477] = 8;
razn_h_mem[2478] = 138;
razn_h_mem[2479] = 14;
razn_h_mem[2480] = 144;
razn_h_mem[2481] = 20;
razn_h_mem[2482] = 150;
razn_h_mem[2483] = 26;
razn_h_mem[2484] = 156;
razn_h_mem[2485] = 32;
razn_h_mem[2486] = 162;
razn_h_mem[2487] = 38;
razn_h_mem[2488] = 168;
razn_h_mem[2489] = 44;
razn_h_mem[2490] = 174;
razn_h_mem[2491] = 50;
razn_h_mem[2492] = 180;
razn_h_mem[2493] = 56;
razn_h_mem[2494] = 186;
razn_h_mem[2495] = 62;
razn_h_mem[2496] = 192;
razn_h_mem[2497] = 68;
razn_h_mem[2498] = 198;
razn_h_mem[2499] = 74;
razn_h_mem[2500] = 204;
razn_h_mem[2501] = 80;
razn_h_mem[2502] = 210;
razn_h_mem[2503] = 86;
razn_h_mem[2504] = 216;
razn_h_mem[2505] = 92;
razn_h_mem[2506] = 222;
razn_h_mem[2507] = 98;
razn_h_mem[2508] = 228;
razn_h_mem[2509] = 104;
razn_h_mem[2510] = 234;
razn_h_mem[2511] = 110;
razn_h_mem[2512] = 240;
razn_h_mem[2513] = 116;
razn_h_mem[2514] = 246;
razn_h_mem[2515] = 122;
razn_h_mem[2516] = 252;
razn_h_mem[2517] = 128;
razn_h_mem[2518] = 4;
razn_h_mem[2519] = 134;
razn_h_mem[2520] = 10;
razn_h_mem[2521] = 140;
razn_h_mem[2522] = 16;
razn_h_mem[2523] = 146;
razn_h_mem[2524] = 22;
razn_h_mem[2525] = 152;
razn_h_mem[2526] = 28;
razn_h_mem[2527] = 158;
razn_h_mem[2528] = 34;
razn_h_mem[2529] = 164;
razn_h_mem[2530] = 40;
razn_h_mem[2531] = 170;
razn_h_mem[2532] = 46;
razn_h_mem[2533] = 176;
razn_h_mem[2534] = 52;
razn_h_mem[2535] = 182;
razn_h_mem[2536] = 58;
razn_h_mem[2537] = 188;
razn_h_mem[2538] = 64;
razn_h_mem[2539] = 194;
razn_h_mem[2540] = 70;
razn_h_mem[2541] = 200;
razn_h_mem[2542] = 76;
razn_h_mem[2543] = 206;
razn_h_mem[2544] = 82;
razn_h_mem[2545] = 212;
razn_h_mem[2546] = 88;
razn_h_mem[2547] = 218;
razn_h_mem[2548] = 94;
razn_h_mem[2549] = 224;
razn_h_mem[2550] = 100;
razn_h_mem[2551] = 230;
razn_h_mem[2552] = 106;
razn_h_mem[2553] = 236;
razn_h_mem[2554] = 112;
razn_h_mem[2555] = 242;
razn_h_mem[2556] = 118;
razn_h_mem[2557] = 248;
razn_h_mem[2558] = 124;
razn_h_mem[2559] = 255;
razn_h_mem[2560] = 0;
razn_h_mem[2561] = 130;
razn_h_mem[2562] = 6;
razn_h_mem[2563] = 136;
razn_h_mem[2564] = 12;
razn_h_mem[2565] = 142;
razn_h_mem[2566] = 18;
razn_h_mem[2567] = 148;
razn_h_mem[2568] = 24;
razn_h_mem[2569] = 154;
razn_h_mem[2570] = 30;
razn_h_mem[2571] = 160;
razn_h_mem[2572] = 36;
razn_h_mem[2573] = 166;
razn_h_mem[2574] = 42;
razn_h_mem[2575] = 172;
razn_h_mem[2576] = 48;
razn_h_mem[2577] = 178;
razn_h_mem[2578] = 54;
razn_h_mem[2579] = 184;
razn_h_mem[2580] = 60;
razn_h_mem[2581] = 190;
razn_h_mem[2582] = 66;
razn_h_mem[2583] = 196;
razn_h_mem[2584] = 72;
razn_h_mem[2585] = 202;
razn_h_mem[2586] = 78;
razn_h_mem[2587] = 208;
razn_h_mem[2588] = 84;
razn_h_mem[2589] = 214;
razn_h_mem[2590] = 90;
razn_h_mem[2591] = 220;
razn_h_mem[2592] = 96;
razn_h_mem[2593] = 226;
razn_h_mem[2594] = 102;
razn_h_mem[2595] = 232;
razn_h_mem[2596] = 108;
razn_h_mem[2597] = 238;
razn_h_mem[2598] = 114;
razn_h_mem[2599] = 244;
razn_h_mem[2600] = 120;
razn_h_mem[2601] = 250;
razn_h_mem[2602] = 126;
razn_h_mem[2603] = 2;
razn_h_mem[2604] = 132;
razn_h_mem[2605] = 8;
razn_h_mem[2606] = 138;
razn_h_mem[2607] = 14;
razn_h_mem[2608] = 144;
razn_h_mem[2609] = 20;
razn_h_mem[2610] = 150;
razn_h_mem[2611] = 26;
razn_h_mem[2612] = 156;
razn_h_mem[2613] = 32;
razn_h_mem[2614] = 162;
razn_h_mem[2615] = 38;
razn_h_mem[2616] = 168;
razn_h_mem[2617] = 44;
razn_h_mem[2618] = 174;
razn_h_mem[2619] = 50;
razn_h_mem[2620] = 180;
razn_h_mem[2621] = 56;
razn_h_mem[2622] = 186;
razn_h_mem[2623] = 62;
razn_h_mem[2624] = 192;
razn_h_mem[2625] = 68;
razn_h_mem[2626] = 198;
razn_h_mem[2627] = 74;
razn_h_mem[2628] = 204;
razn_h_mem[2629] = 80;
razn_h_mem[2630] = 210;
razn_h_mem[2631] = 86;
razn_h_mem[2632] = 216;
razn_h_mem[2633] = 92;
razn_h_mem[2634] = 222;
razn_h_mem[2635] = 98;
razn_h_mem[2636] = 228;
razn_h_mem[2637] = 104;
razn_h_mem[2638] = 234;
razn_h_mem[2639] = 110;
razn_h_mem[2640] = 240;
razn_h_mem[2641] = 116;
razn_h_mem[2642] = 246;
razn_h_mem[2643] = 122;
razn_h_mem[2644] = 252;
razn_h_mem[2645] = 128;
razn_h_mem[2646] = 4;
razn_h_mem[2647] = 134;
razn_h_mem[2648] = 10;
razn_h_mem[2649] = 140;
razn_h_mem[2650] = 16;
razn_h_mem[2651] = 146;
razn_h_mem[2652] = 22;
razn_h_mem[2653] = 152;
razn_h_mem[2654] = 28;
razn_h_mem[2655] = 158;
razn_h_mem[2656] = 34;
razn_h_mem[2657] = 164;
razn_h_mem[2658] = 40;
razn_h_mem[2659] = 170;
razn_h_mem[2660] = 46;
razn_h_mem[2661] = 176;
razn_h_mem[2662] = 52;
razn_h_mem[2663] = 182;
razn_h_mem[2664] = 58;
razn_h_mem[2665] = 188;
razn_h_mem[2666] = 64;
razn_h_mem[2667] = 194;
razn_h_mem[2668] = 70;
razn_h_mem[2669] = 200;
razn_h_mem[2670] = 76;
razn_h_mem[2671] = 206;
razn_h_mem[2672] = 82;
razn_h_mem[2673] = 212;
razn_h_mem[2674] = 88;
razn_h_mem[2675] = 218;
razn_h_mem[2676] = 94;
razn_h_mem[2677] = 224;
razn_h_mem[2678] = 100;
razn_h_mem[2679] = 230;
razn_h_mem[2680] = 106;
razn_h_mem[2681] = 236;
razn_h_mem[2682] = 112;
razn_h_mem[2683] = 242;
razn_h_mem[2684] = 118;
razn_h_mem[2685] = 248;
razn_h_mem[2686] = 124;
razn_h_mem[2687] = 255;
razn_h_mem[2688] = 0;
razn_h_mem[2689] = 130;
razn_h_mem[2690] = 6;
razn_h_mem[2691] = 136;
razn_h_mem[2692] = 12;
razn_h_mem[2693] = 142;
razn_h_mem[2694] = 18;
razn_h_mem[2695] = 148;
razn_h_mem[2696] = 24;
razn_h_mem[2697] = 154;
razn_h_mem[2698] = 30;
razn_h_mem[2699] = 160;
razn_h_mem[2700] = 36;
razn_h_mem[2701] = 166;
razn_h_mem[2702] = 42;
razn_h_mem[2703] = 172;
razn_h_mem[2704] = 48;
razn_h_mem[2705] = 178;
razn_h_mem[2706] = 54;
razn_h_mem[2707] = 184;
razn_h_mem[2708] = 60;
razn_h_mem[2709] = 190;
razn_h_mem[2710] = 66;
razn_h_mem[2711] = 196;
razn_h_mem[2712] = 72;
razn_h_mem[2713] = 202;
razn_h_mem[2714] = 78;
razn_h_mem[2715] = 208;
razn_h_mem[2716] = 84;
razn_h_mem[2717] = 214;
razn_h_mem[2718] = 90;
razn_h_mem[2719] = 220;
razn_h_mem[2720] = 96;
razn_h_mem[2721] = 226;
razn_h_mem[2722] = 102;
razn_h_mem[2723] = 232;
razn_h_mem[2724] = 108;
razn_h_mem[2725] = 238;
razn_h_mem[2726] = 114;
razn_h_mem[2727] = 244;
razn_h_mem[2728] = 120;
razn_h_mem[2729] = 250;
razn_h_mem[2730] = 126;
razn_h_mem[2731] = 2;
razn_h_mem[2732] = 132;
razn_h_mem[2733] = 8;
razn_h_mem[2734] = 138;
razn_h_mem[2735] = 14;
razn_h_mem[2736] = 144;
razn_h_mem[2737] = 20;
razn_h_mem[2738] = 150;
razn_h_mem[2739] = 26;
razn_h_mem[2740] = 156;
razn_h_mem[2741] = 32;
razn_h_mem[2742] = 162;
razn_h_mem[2743] = 38;
razn_h_mem[2744] = 168;
razn_h_mem[2745] = 44;
razn_h_mem[2746] = 174;
razn_h_mem[2747] = 50;
razn_h_mem[2748] = 180;
razn_h_mem[2749] = 56;
razn_h_mem[2750] = 186;
razn_h_mem[2751] = 62;
razn_h_mem[2752] = 192;
razn_h_mem[2753] = 68;
razn_h_mem[2754] = 198;
razn_h_mem[2755] = 74;
razn_h_mem[2756] = 204;
razn_h_mem[2757] = 80;
razn_h_mem[2758] = 210;
razn_h_mem[2759] = 86;
razn_h_mem[2760] = 216;
razn_h_mem[2761] = 92;
razn_h_mem[2762] = 222;
razn_h_mem[2763] = 98;
razn_h_mem[2764] = 228;
razn_h_mem[2765] = 104;
razn_h_mem[2766] = 234;
razn_h_mem[2767] = 110;
razn_h_mem[2768] = 240;
razn_h_mem[2769] = 116;
razn_h_mem[2770] = 246;
razn_h_mem[2771] = 122;
razn_h_mem[2772] = 252;
razn_h_mem[2773] = 128;
razn_h_mem[2774] = 4;
razn_h_mem[2775] = 134;
razn_h_mem[2776] = 10;
razn_h_mem[2777] = 140;
razn_h_mem[2778] = 16;
razn_h_mem[2779] = 146;
razn_h_mem[2780] = 22;
razn_h_mem[2781] = 152;
razn_h_mem[2782] = 28;
razn_h_mem[2783] = 158;
razn_h_mem[2784] = 34;
razn_h_mem[2785] = 164;
razn_h_mem[2786] = 40;
razn_h_mem[2787] = 170;
razn_h_mem[2788] = 46;
razn_h_mem[2789] = 176;
razn_h_mem[2790] = 52;
razn_h_mem[2791] = 182;
razn_h_mem[2792] = 58;
razn_h_mem[2793] = 188;
razn_h_mem[2794] = 64;
razn_h_mem[2795] = 194;
razn_h_mem[2796] = 70;
razn_h_mem[2797] = 200;
razn_h_mem[2798] = 76;
razn_h_mem[2799] = 206;
razn_h_mem[2800] = 82;
razn_h_mem[2801] = 212;
razn_h_mem[2802] = 88;
razn_h_mem[2803] = 218;
razn_h_mem[2804] = 94;
razn_h_mem[2805] = 224;
razn_h_mem[2806] = 100;
razn_h_mem[2807] = 230;
razn_h_mem[2808] = 106;
razn_h_mem[2809] = 236;
razn_h_mem[2810] = 112;
razn_h_mem[2811] = 242;
razn_h_mem[2812] = 118;
razn_h_mem[2813] = 248;
razn_h_mem[2814] = 124;
razn_h_mem[2815] = 255;
razn_h_mem[2816] = 0;
razn_h_mem[2817] = 130;
razn_h_mem[2818] = 6;
razn_h_mem[2819] = 136;
razn_h_mem[2820] = 12;
razn_h_mem[2821] = 142;
razn_h_mem[2822] = 18;
razn_h_mem[2823] = 148;
razn_h_mem[2824] = 24;
razn_h_mem[2825] = 154;
razn_h_mem[2826] = 30;
razn_h_mem[2827] = 160;
razn_h_mem[2828] = 36;
razn_h_mem[2829] = 166;
razn_h_mem[2830] = 42;
razn_h_mem[2831] = 172;
razn_h_mem[2832] = 48;
razn_h_mem[2833] = 178;
razn_h_mem[2834] = 54;
razn_h_mem[2835] = 184;
razn_h_mem[2836] = 60;
razn_h_mem[2837] = 190;
razn_h_mem[2838] = 66;
razn_h_mem[2839] = 196;
razn_h_mem[2840] = 72;
razn_h_mem[2841] = 202;
razn_h_mem[2842] = 78;
razn_h_mem[2843] = 208;
razn_h_mem[2844] = 84;
razn_h_mem[2845] = 214;
razn_h_mem[2846] = 90;
razn_h_mem[2847] = 220;
razn_h_mem[2848] = 96;
razn_h_mem[2849] = 226;
razn_h_mem[2850] = 102;
razn_h_mem[2851] = 232;
razn_h_mem[2852] = 108;
razn_h_mem[2853] = 238;
razn_h_mem[2854] = 114;
razn_h_mem[2855] = 244;
razn_h_mem[2856] = 120;
razn_h_mem[2857] = 250;
razn_h_mem[2858] = 126;
razn_h_mem[2859] = 2;
razn_h_mem[2860] = 132;
razn_h_mem[2861] = 8;
razn_h_mem[2862] = 138;
razn_h_mem[2863] = 14;
razn_h_mem[2864] = 144;
razn_h_mem[2865] = 20;
razn_h_mem[2866] = 150;
razn_h_mem[2867] = 26;
razn_h_mem[2868] = 156;
razn_h_mem[2869] = 32;
razn_h_mem[2870] = 162;
razn_h_mem[2871] = 38;
razn_h_mem[2872] = 168;
razn_h_mem[2873] = 44;
razn_h_mem[2874] = 174;
razn_h_mem[2875] = 50;
razn_h_mem[2876] = 180;
razn_h_mem[2877] = 56;
razn_h_mem[2878] = 186;
razn_h_mem[2879] = 62;
razn_h_mem[2880] = 192;
razn_h_mem[2881] = 68;
razn_h_mem[2882] = 198;
razn_h_mem[2883] = 74;
razn_h_mem[2884] = 204;
razn_h_mem[2885] = 80;
razn_h_mem[2886] = 210;
razn_h_mem[2887] = 86;
razn_h_mem[2888] = 216;
razn_h_mem[2889] = 92;
razn_h_mem[2890] = 222;
razn_h_mem[2891] = 98;
razn_h_mem[2892] = 228;
razn_h_mem[2893] = 104;
razn_h_mem[2894] = 234;
razn_h_mem[2895] = 110;
razn_h_mem[2896] = 240;
razn_h_mem[2897] = 116;
razn_h_mem[2898] = 246;
razn_h_mem[2899] = 122;
razn_h_mem[2900] = 252;
razn_h_mem[2901] = 128;
razn_h_mem[2902] = 4;
razn_h_mem[2903] = 134;
razn_h_mem[2904] = 10;
razn_h_mem[2905] = 140;
razn_h_mem[2906] = 16;
razn_h_mem[2907] = 146;
razn_h_mem[2908] = 22;
razn_h_mem[2909] = 152;
razn_h_mem[2910] = 28;
razn_h_mem[2911] = 158;
razn_h_mem[2912] = 34;
razn_h_mem[2913] = 164;
razn_h_mem[2914] = 40;
razn_h_mem[2915] = 170;
razn_h_mem[2916] = 46;
razn_h_mem[2917] = 176;
razn_h_mem[2918] = 52;
razn_h_mem[2919] = 182;
razn_h_mem[2920] = 58;
razn_h_mem[2921] = 188;
razn_h_mem[2922] = 64;
razn_h_mem[2923] = 194;
razn_h_mem[2924] = 70;
razn_h_mem[2925] = 200;
razn_h_mem[2926] = 76;
razn_h_mem[2927] = 206;
razn_h_mem[2928] = 82;
razn_h_mem[2929] = 212;
razn_h_mem[2930] = 88;
razn_h_mem[2931] = 218;
razn_h_mem[2932] = 94;
razn_h_mem[2933] = 224;
razn_h_mem[2934] = 100;
razn_h_mem[2935] = 230;
razn_h_mem[2936] = 106;
razn_h_mem[2937] = 236;
razn_h_mem[2938] = 112;
razn_h_mem[2939] = 242;
razn_h_mem[2940] = 118;
razn_h_mem[2941] = 248;
razn_h_mem[2942] = 124;
razn_h_mem[2943] = 255;
razn_h_mem[2944] = 0;
razn_h_mem[2945] = 130;
razn_h_mem[2946] = 6;
razn_h_mem[2947] = 136;
razn_h_mem[2948] = 12;
razn_h_mem[2949] = 142;
razn_h_mem[2950] = 18;
razn_h_mem[2951] = 148;
razn_h_mem[2952] = 24;
razn_h_mem[2953] = 154;
razn_h_mem[2954] = 30;
razn_h_mem[2955] = 160;
razn_h_mem[2956] = 36;
razn_h_mem[2957] = 166;
razn_h_mem[2958] = 42;
razn_h_mem[2959] = 172;
razn_h_mem[2960] = 48;
razn_h_mem[2961] = 178;
razn_h_mem[2962] = 54;
razn_h_mem[2963] = 184;
razn_h_mem[2964] = 60;
razn_h_mem[2965] = 190;
razn_h_mem[2966] = 66;
razn_h_mem[2967] = 196;
razn_h_mem[2968] = 72;
razn_h_mem[2969] = 202;
razn_h_mem[2970] = 78;
razn_h_mem[2971] = 208;
razn_h_mem[2972] = 84;
razn_h_mem[2973] = 214;
razn_h_mem[2974] = 90;
razn_h_mem[2975] = 220;
razn_h_mem[2976] = 96;
razn_h_mem[2977] = 226;
razn_h_mem[2978] = 102;
razn_h_mem[2979] = 232;
razn_h_mem[2980] = 108;
razn_h_mem[2981] = 238;
razn_h_mem[2982] = 114;
razn_h_mem[2983] = 244;
razn_h_mem[2984] = 120;
razn_h_mem[2985] = 250;
razn_h_mem[2986] = 126;
razn_h_mem[2987] = 2;
razn_h_mem[2988] = 132;
razn_h_mem[2989] = 8;
razn_h_mem[2990] = 138;
razn_h_mem[2991] = 14;
razn_h_mem[2992] = 144;
razn_h_mem[2993] = 20;
razn_h_mem[2994] = 150;
razn_h_mem[2995] = 26;
razn_h_mem[2996] = 156;
razn_h_mem[2997] = 32;
razn_h_mem[2998] = 162;
razn_h_mem[2999] = 38;
razn_h_mem[3000] = 168;
razn_h_mem[3001] = 44;
razn_h_mem[3002] = 174;
razn_h_mem[3003] = 50;
razn_h_mem[3004] = 180;
razn_h_mem[3005] = 56;
razn_h_mem[3006] = 186;
razn_h_mem[3007] = 62;
razn_h_mem[3008] = 192;
razn_h_mem[3009] = 68;
razn_h_mem[3010] = 198;
razn_h_mem[3011] = 74;
razn_h_mem[3012] = 204;
razn_h_mem[3013] = 80;
razn_h_mem[3014] = 210;
razn_h_mem[3015] = 86;
razn_h_mem[3016] = 216;
razn_h_mem[3017] = 92;
razn_h_mem[3018] = 222;
razn_h_mem[3019] = 98;
razn_h_mem[3020] = 228;
razn_h_mem[3021] = 104;
razn_h_mem[3022] = 234;
razn_h_mem[3023] = 110;
razn_h_mem[3024] = 240;
razn_h_mem[3025] = 116;
razn_h_mem[3026] = 246;
razn_h_mem[3027] = 122;
razn_h_mem[3028] = 252;
razn_h_mem[3029] = 128;
razn_h_mem[3030] = 4;
razn_h_mem[3031] = 134;
razn_h_mem[3032] = 10;
razn_h_mem[3033] = 140;
razn_h_mem[3034] = 16;
razn_h_mem[3035] = 146;
razn_h_mem[3036] = 22;
razn_h_mem[3037] = 152;
razn_h_mem[3038] = 28;
razn_h_mem[3039] = 158;
razn_h_mem[3040] = 34;
razn_h_mem[3041] = 164;
razn_h_mem[3042] = 40;
razn_h_mem[3043] = 170;
razn_h_mem[3044] = 46;
razn_h_mem[3045] = 176;
razn_h_mem[3046] = 52;
razn_h_mem[3047] = 182;
razn_h_mem[3048] = 58;
razn_h_mem[3049] = 188;
razn_h_mem[3050] = 64;
razn_h_mem[3051] = 194;
razn_h_mem[3052] = 70;
razn_h_mem[3053] = 200;
razn_h_mem[3054] = 76;
razn_h_mem[3055] = 206;
razn_h_mem[3056] = 82;
razn_h_mem[3057] = 212;
razn_h_mem[3058] = 88;
razn_h_mem[3059] = 218;
razn_h_mem[3060] = 94;
razn_h_mem[3061] = 224;
razn_h_mem[3062] = 100;
razn_h_mem[3063] = 230;
razn_h_mem[3064] = 106;
razn_h_mem[3065] = 236;
razn_h_mem[3066] = 112;
razn_h_mem[3067] = 242;
razn_h_mem[3068] = 118;
razn_h_mem[3069] = 248;
razn_h_mem[3070] = 124;
razn_h_mem[3071] = 255;
razn_h_mem[3072] = 0;
razn_h_mem[3073] = 130;
razn_h_mem[3074] = 6;
razn_h_mem[3075] = 136;
razn_h_mem[3076] = 12;
razn_h_mem[3077] = 142;
razn_h_mem[3078] = 18;
razn_h_mem[3079] = 148;
razn_h_mem[3080] = 24;
razn_h_mem[3081] = 154;
razn_h_mem[3082] = 30;
razn_h_mem[3083] = 160;
razn_h_mem[3084] = 36;
razn_h_mem[3085] = 166;
razn_h_mem[3086] = 42;
razn_h_mem[3087] = 172;
razn_h_mem[3088] = 48;
razn_h_mem[3089] = 178;
razn_h_mem[3090] = 54;
razn_h_mem[3091] = 184;
razn_h_mem[3092] = 60;
razn_h_mem[3093] = 190;
razn_h_mem[3094] = 66;
razn_h_mem[3095] = 196;
razn_h_mem[3096] = 72;
razn_h_mem[3097] = 202;
razn_h_mem[3098] = 78;
razn_h_mem[3099] = 208;
razn_h_mem[3100] = 84;
razn_h_mem[3101] = 214;
razn_h_mem[3102] = 90;
razn_h_mem[3103] = 220;
razn_h_mem[3104] = 96;
razn_h_mem[3105] = 226;
razn_h_mem[3106] = 102;
razn_h_mem[3107] = 232;
razn_h_mem[3108] = 108;
razn_h_mem[3109] = 238;
razn_h_mem[3110] = 114;
razn_h_mem[3111] = 244;
razn_h_mem[3112] = 120;
razn_h_mem[3113] = 250;
razn_h_mem[3114] = 126;
razn_h_mem[3115] = 2;
razn_h_mem[3116] = 132;
razn_h_mem[3117] = 8;
razn_h_mem[3118] = 138;
razn_h_mem[3119] = 14;
razn_h_mem[3120] = 144;
razn_h_mem[3121] = 20;
razn_h_mem[3122] = 150;
razn_h_mem[3123] = 26;
razn_h_mem[3124] = 156;
razn_h_mem[3125] = 32;
razn_h_mem[3126] = 162;
razn_h_mem[3127] = 38;
razn_h_mem[3128] = 168;
razn_h_mem[3129] = 44;
razn_h_mem[3130] = 174;
razn_h_mem[3131] = 50;
razn_h_mem[3132] = 180;
razn_h_mem[3133] = 56;
razn_h_mem[3134] = 186;
razn_h_mem[3135] = 62;
razn_h_mem[3136] = 192;
razn_h_mem[3137] = 68;
razn_h_mem[3138] = 198;
razn_h_mem[3139] = 74;
razn_h_mem[3140] = 204;
razn_h_mem[3141] = 80;
razn_h_mem[3142] = 210;
razn_h_mem[3143] = 86;
razn_h_mem[3144] = 216;
razn_h_mem[3145] = 92;
razn_h_mem[3146] = 222;
razn_h_mem[3147] = 98;
razn_h_mem[3148] = 228;
razn_h_mem[3149] = 104;
razn_h_mem[3150] = 234;
razn_h_mem[3151] = 110;
razn_h_mem[3152] = 240;
razn_h_mem[3153] = 116;
razn_h_mem[3154] = 246;
razn_h_mem[3155] = 122;
razn_h_mem[3156] = 252;
razn_h_mem[3157] = 128;
razn_h_mem[3158] = 4;
razn_h_mem[3159] = 134;
razn_h_mem[3160] = 10;
razn_h_mem[3161] = 140;
razn_h_mem[3162] = 16;
razn_h_mem[3163] = 146;
razn_h_mem[3164] = 22;
razn_h_mem[3165] = 152;
razn_h_mem[3166] = 28;
razn_h_mem[3167] = 158;
razn_h_mem[3168] = 34;
razn_h_mem[3169] = 164;
razn_h_mem[3170] = 40;
razn_h_mem[3171] = 170;
razn_h_mem[3172] = 46;
razn_h_mem[3173] = 176;
razn_h_mem[3174] = 52;
razn_h_mem[3175] = 182;
razn_h_mem[3176] = 58;
razn_h_mem[3177] = 188;
razn_h_mem[3178] = 64;
razn_h_mem[3179] = 194;
razn_h_mem[3180] = 70;
razn_h_mem[3181] = 200;
razn_h_mem[3182] = 76;
razn_h_mem[3183] = 206;
razn_h_mem[3184] = 82;
razn_h_mem[3185] = 212;
razn_h_mem[3186] = 88;
razn_h_mem[3187] = 218;
razn_h_mem[3188] = 94;
razn_h_mem[3189] = 224;
razn_h_mem[3190] = 100;
razn_h_mem[3191] = 230;
razn_h_mem[3192] = 106;
razn_h_mem[3193] = 236;
razn_h_mem[3194] = 112;
razn_h_mem[3195] = 242;
razn_h_mem[3196] = 118;
razn_h_mem[3197] = 248;
razn_h_mem[3198] = 124;
razn_h_mem[3199] = 255;
razn_h_mem[3200] = 0;
razn_h_mem[3201] = 130;
razn_h_mem[3202] = 6;
razn_h_mem[3203] = 136;
razn_h_mem[3204] = 12;
razn_h_mem[3205] = 142;
razn_h_mem[3206] = 18;
razn_h_mem[3207] = 148;
razn_h_mem[3208] = 24;
razn_h_mem[3209] = 154;
razn_h_mem[3210] = 30;
razn_h_mem[3211] = 160;
razn_h_mem[3212] = 36;
razn_h_mem[3213] = 166;
razn_h_mem[3214] = 42;
razn_h_mem[3215] = 172;
razn_h_mem[3216] = 48;
razn_h_mem[3217] = 178;
razn_h_mem[3218] = 54;
razn_h_mem[3219] = 184;
razn_h_mem[3220] = 60;
razn_h_mem[3221] = 190;
razn_h_mem[3222] = 66;
razn_h_mem[3223] = 196;
razn_h_mem[3224] = 72;
razn_h_mem[3225] = 202;
razn_h_mem[3226] = 78;
razn_h_mem[3227] = 208;
razn_h_mem[3228] = 84;
razn_h_mem[3229] = 214;
razn_h_mem[3230] = 90;
razn_h_mem[3231] = 220;
razn_h_mem[3232] = 96;
razn_h_mem[3233] = 226;
razn_h_mem[3234] = 102;
razn_h_mem[3235] = 232;
razn_h_mem[3236] = 108;
razn_h_mem[3237] = 238;
razn_h_mem[3238] = 114;
razn_h_mem[3239] = 244;
razn_h_mem[3240] = 120;
razn_h_mem[3241] = 250;
razn_h_mem[3242] = 126;
razn_h_mem[3243] = 2;
razn_h_mem[3244] = 132;
razn_h_mem[3245] = 8;
razn_h_mem[3246] = 138;
razn_h_mem[3247] = 14;
razn_h_mem[3248] = 144;
razn_h_mem[3249] = 20;
razn_h_mem[3250] = 150;
razn_h_mem[3251] = 26;
razn_h_mem[3252] = 156;
razn_h_mem[3253] = 32;
razn_h_mem[3254] = 162;
razn_h_mem[3255] = 38;
razn_h_mem[3256] = 168;
razn_h_mem[3257] = 44;
razn_h_mem[3258] = 174;
razn_h_mem[3259] = 50;
razn_h_mem[3260] = 180;
razn_h_mem[3261] = 56;
razn_h_mem[3262] = 186;
razn_h_mem[3263] = 62;
razn_h_mem[3264] = 192;
razn_h_mem[3265] = 68;
razn_h_mem[3266] = 198;
razn_h_mem[3267] = 74;
razn_h_mem[3268] = 204;
razn_h_mem[3269] = 80;
razn_h_mem[3270] = 210;
razn_h_mem[3271] = 86;
razn_h_mem[3272] = 216;
razn_h_mem[3273] = 92;
razn_h_mem[3274] = 222;
razn_h_mem[3275] = 98;
razn_h_mem[3276] = 228;
razn_h_mem[3277] = 104;
razn_h_mem[3278] = 234;
razn_h_mem[3279] = 110;
razn_h_mem[3280] = 240;
razn_h_mem[3281] = 116;
razn_h_mem[3282] = 246;
razn_h_mem[3283] = 122;
razn_h_mem[3284] = 252;
razn_h_mem[3285] = 128;
razn_h_mem[3286] = 4;
razn_h_mem[3287] = 134;
razn_h_mem[3288] = 10;
razn_h_mem[3289] = 140;
razn_h_mem[3290] = 16;
razn_h_mem[3291] = 146;
razn_h_mem[3292] = 22;
razn_h_mem[3293] = 152;
razn_h_mem[3294] = 28;
razn_h_mem[3295] = 158;
razn_h_mem[3296] = 34;
razn_h_mem[3297] = 164;
razn_h_mem[3298] = 40;
razn_h_mem[3299] = 170;
razn_h_mem[3300] = 46;
razn_h_mem[3301] = 176;
razn_h_mem[3302] = 52;
razn_h_mem[3303] = 182;
razn_h_mem[3304] = 58;
razn_h_mem[3305] = 188;
razn_h_mem[3306] = 64;
razn_h_mem[3307] = 194;
razn_h_mem[3308] = 70;
razn_h_mem[3309] = 200;
razn_h_mem[3310] = 76;
razn_h_mem[3311] = 206;
razn_h_mem[3312] = 82;
razn_h_mem[3313] = 212;
razn_h_mem[3314] = 88;
razn_h_mem[3315] = 218;
razn_h_mem[3316] = 94;
razn_h_mem[3317] = 224;
razn_h_mem[3318] = 100;
razn_h_mem[3319] = 230;
razn_h_mem[3320] = 106;
razn_h_mem[3321] = 236;
razn_h_mem[3322] = 112;
razn_h_mem[3323] = 242;
razn_h_mem[3324] = 118;
razn_h_mem[3325] = 248;
razn_h_mem[3326] = 124;
razn_h_mem[3327] = 255;
razn_h_mem[3328] = 0;
razn_h_mem[3329] = 130;
razn_h_mem[3330] = 6;
razn_h_mem[3331] = 136;
razn_h_mem[3332] = 12;
razn_h_mem[3333] = 142;
razn_h_mem[3334] = 18;
razn_h_mem[3335] = 148;
razn_h_mem[3336] = 24;
razn_h_mem[3337] = 154;
razn_h_mem[3338] = 30;
razn_h_mem[3339] = 160;
razn_h_mem[3340] = 36;
razn_h_mem[3341] = 166;
razn_h_mem[3342] = 42;
razn_h_mem[3343] = 172;
razn_h_mem[3344] = 48;
razn_h_mem[3345] = 178;
razn_h_mem[3346] = 54;
razn_h_mem[3347] = 184;
razn_h_mem[3348] = 60;
razn_h_mem[3349] = 190;
razn_h_mem[3350] = 66;
razn_h_mem[3351] = 196;
razn_h_mem[3352] = 72;
razn_h_mem[3353] = 202;
razn_h_mem[3354] = 78;
razn_h_mem[3355] = 208;
razn_h_mem[3356] = 84;
razn_h_mem[3357] = 214;
razn_h_mem[3358] = 90;
razn_h_mem[3359] = 220;
razn_h_mem[3360] = 96;
razn_h_mem[3361] = 226;
razn_h_mem[3362] = 102;
razn_h_mem[3363] = 232;
razn_h_mem[3364] = 108;
razn_h_mem[3365] = 238;
razn_h_mem[3366] = 114;
razn_h_mem[3367] = 244;
razn_h_mem[3368] = 120;
razn_h_mem[3369] = 250;
razn_h_mem[3370] = 126;
razn_h_mem[3371] = 2;
razn_h_mem[3372] = 132;
razn_h_mem[3373] = 8;
razn_h_mem[3374] = 138;
razn_h_mem[3375] = 14;
razn_h_mem[3376] = 144;
razn_h_mem[3377] = 20;
razn_h_mem[3378] = 150;
razn_h_mem[3379] = 26;
razn_h_mem[3380] = 156;
razn_h_mem[3381] = 32;
razn_h_mem[3382] = 162;
razn_h_mem[3383] = 38;
razn_h_mem[3384] = 168;
razn_h_mem[3385] = 44;
razn_h_mem[3386] = 174;
razn_h_mem[3387] = 50;
razn_h_mem[3388] = 180;
razn_h_mem[3389] = 56;
razn_h_mem[3390] = 186;
razn_h_mem[3391] = 62;
razn_h_mem[3392] = 192;
razn_h_mem[3393] = 68;
razn_h_mem[3394] = 198;
razn_h_mem[3395] = 74;
razn_h_mem[3396] = 204;
razn_h_mem[3397] = 80;
razn_h_mem[3398] = 210;
razn_h_mem[3399] = 86;
razn_h_mem[3400] = 216;
razn_h_mem[3401] = 92;
razn_h_mem[3402] = 222;
razn_h_mem[3403] = 98;
razn_h_mem[3404] = 228;
razn_h_mem[3405] = 104;
razn_h_mem[3406] = 234;
razn_h_mem[3407] = 110;
razn_h_mem[3408] = 240;
razn_h_mem[3409] = 116;
razn_h_mem[3410] = 246;
razn_h_mem[3411] = 122;
razn_h_mem[3412] = 252;
razn_h_mem[3413] = 128;
razn_h_mem[3414] = 4;
razn_h_mem[3415] = 134;
razn_h_mem[3416] = 10;
razn_h_mem[3417] = 140;
razn_h_mem[3418] = 16;
razn_h_mem[3419] = 146;
razn_h_mem[3420] = 22;
razn_h_mem[3421] = 152;
razn_h_mem[3422] = 28;
razn_h_mem[3423] = 158;
razn_h_mem[3424] = 34;
razn_h_mem[3425] = 164;
razn_h_mem[3426] = 40;
razn_h_mem[3427] = 170;
razn_h_mem[3428] = 46;
razn_h_mem[3429] = 176;
razn_h_mem[3430] = 52;
razn_h_mem[3431] = 182;
razn_h_mem[3432] = 58;
razn_h_mem[3433] = 188;
razn_h_mem[3434] = 64;
razn_h_mem[3435] = 194;
razn_h_mem[3436] = 70;
razn_h_mem[3437] = 200;
razn_h_mem[3438] = 76;
razn_h_mem[3439] = 206;
razn_h_mem[3440] = 82;
razn_h_mem[3441] = 212;
razn_h_mem[3442] = 88;
razn_h_mem[3443] = 218;
razn_h_mem[3444] = 94;
razn_h_mem[3445] = 224;
razn_h_mem[3446] = 100;
razn_h_mem[3447] = 230;
razn_h_mem[3448] = 106;
razn_h_mem[3449] = 236;
razn_h_mem[3450] = 112;
razn_h_mem[3451] = 242;
razn_h_mem[3452] = 118;
razn_h_mem[3453] = 248;
razn_h_mem[3454] = 124;
razn_h_mem[3455] = 255;
razn_h_mem[3456] = 0;
razn_h_mem[3457] = 130;
razn_h_mem[3458] = 6;
razn_h_mem[3459] = 136;
razn_h_mem[3460] = 12;
razn_h_mem[3461] = 142;
razn_h_mem[3462] = 18;
razn_h_mem[3463] = 148;
razn_h_mem[3464] = 24;
razn_h_mem[3465] = 154;
razn_h_mem[3466] = 30;
razn_h_mem[3467] = 160;
razn_h_mem[3468] = 36;
razn_h_mem[3469] = 166;
razn_h_mem[3470] = 42;
razn_h_mem[3471] = 172;
razn_h_mem[3472] = 48;
razn_h_mem[3473] = 178;
razn_h_mem[3474] = 54;
razn_h_mem[3475] = 184;
razn_h_mem[3476] = 60;
razn_h_mem[3477] = 190;
razn_h_mem[3478] = 66;
razn_h_mem[3479] = 196;
razn_h_mem[3480] = 72;
razn_h_mem[3481] = 202;
razn_h_mem[3482] = 78;
razn_h_mem[3483] = 208;
razn_h_mem[3484] = 84;
razn_h_mem[3485] = 214;
razn_h_mem[3486] = 90;
razn_h_mem[3487] = 220;
razn_h_mem[3488] = 96;
razn_h_mem[3489] = 226;
razn_h_mem[3490] = 102;
razn_h_mem[3491] = 232;
razn_h_mem[3492] = 108;
razn_h_mem[3493] = 238;
razn_h_mem[3494] = 114;
razn_h_mem[3495] = 244;
razn_h_mem[3496] = 120;
razn_h_mem[3497] = 250;
razn_h_mem[3498] = 126;
razn_h_mem[3499] = 2;
razn_h_mem[3500] = 132;
razn_h_mem[3501] = 8;
razn_h_mem[3502] = 138;
razn_h_mem[3503] = 14;
razn_h_mem[3504] = 144;
razn_h_mem[3505] = 20;
razn_h_mem[3506] = 150;
razn_h_mem[3507] = 26;
razn_h_mem[3508] = 156;
razn_h_mem[3509] = 32;
razn_h_mem[3510] = 162;
razn_h_mem[3511] = 38;
razn_h_mem[3512] = 168;
razn_h_mem[3513] = 44;
razn_h_mem[3514] = 174;
razn_h_mem[3515] = 50;
razn_h_mem[3516] = 180;
razn_h_mem[3517] = 56;
razn_h_mem[3518] = 186;
razn_h_mem[3519] = 62;
razn_h_mem[3520] = 192;
razn_h_mem[3521] = 68;
razn_h_mem[3522] = 198;
razn_h_mem[3523] = 74;
razn_h_mem[3524] = 204;
razn_h_mem[3525] = 80;
razn_h_mem[3526] = 210;
razn_h_mem[3527] = 86;
razn_h_mem[3528] = 216;
razn_h_mem[3529] = 92;
razn_h_mem[3530] = 222;
razn_h_mem[3531] = 98;
razn_h_mem[3532] = 228;
razn_h_mem[3533] = 104;
razn_h_mem[3534] = 234;
razn_h_mem[3535] = 110;
razn_h_mem[3536] = 240;
razn_h_mem[3537] = 116;
razn_h_mem[3538] = 246;
razn_h_mem[3539] = 122;
razn_h_mem[3540] = 252;
razn_h_mem[3541] = 128;
razn_h_mem[3542] = 4;
razn_h_mem[3543] = 134;
razn_h_mem[3544] = 10;
razn_h_mem[3545] = 140;
razn_h_mem[3546] = 16;
razn_h_mem[3547] = 146;
razn_h_mem[3548] = 22;
razn_h_mem[3549] = 152;
razn_h_mem[3550] = 28;
razn_h_mem[3551] = 158;
razn_h_mem[3552] = 34;
razn_h_mem[3553] = 164;
razn_h_mem[3554] = 40;
razn_h_mem[3555] = 170;
razn_h_mem[3556] = 46;
razn_h_mem[3557] = 176;
razn_h_mem[3558] = 52;
razn_h_mem[3559] = 182;
razn_h_mem[3560] = 58;
razn_h_mem[3561] = 188;
razn_h_mem[3562] = 64;
razn_h_mem[3563] = 194;
razn_h_mem[3564] = 70;
razn_h_mem[3565] = 200;
razn_h_mem[3566] = 76;
razn_h_mem[3567] = 206;
razn_h_mem[3568] = 82;
razn_h_mem[3569] = 212;
razn_h_mem[3570] = 88;
razn_h_mem[3571] = 218;
razn_h_mem[3572] = 94;
razn_h_mem[3573] = 224;
razn_h_mem[3574] = 100;
razn_h_mem[3575] = 230;
razn_h_mem[3576] = 106;
razn_h_mem[3577] = 236;
razn_h_mem[3578] = 112;
razn_h_mem[3579] = 242;
razn_h_mem[3580] = 118;
razn_h_mem[3581] = 248;
razn_h_mem[3582] = 124;
razn_h_mem[3583] = 255;
razn_h_mem[3584] = 0;
razn_h_mem[3585] = 130;
razn_h_mem[3586] = 6;
razn_h_mem[3587] = 136;
razn_h_mem[3588] = 12;
razn_h_mem[3589] = 142;
razn_h_mem[3590] = 18;
razn_h_mem[3591] = 148;
razn_h_mem[3592] = 24;
razn_h_mem[3593] = 154;
razn_h_mem[3594] = 30;
razn_h_mem[3595] = 160;
razn_h_mem[3596] = 36;
razn_h_mem[3597] = 166;
razn_h_mem[3598] = 42;
razn_h_mem[3599] = 172;
razn_h_mem[3600] = 48;
razn_h_mem[3601] = 178;
razn_h_mem[3602] = 54;
razn_h_mem[3603] = 184;
razn_h_mem[3604] = 60;
razn_h_mem[3605] = 190;
razn_h_mem[3606] = 66;
razn_h_mem[3607] = 196;
razn_h_mem[3608] = 72;
razn_h_mem[3609] = 202;
razn_h_mem[3610] = 78;
razn_h_mem[3611] = 208;
razn_h_mem[3612] = 84;
razn_h_mem[3613] = 214;
razn_h_mem[3614] = 90;
razn_h_mem[3615] = 220;
razn_h_mem[3616] = 96;
razn_h_mem[3617] = 226;
razn_h_mem[3618] = 102;
razn_h_mem[3619] = 232;
razn_h_mem[3620] = 108;
razn_h_mem[3621] = 238;
razn_h_mem[3622] = 114;
razn_h_mem[3623] = 244;
razn_h_mem[3624] = 120;
razn_h_mem[3625] = 250;
razn_h_mem[3626] = 126;
razn_h_mem[3627] = 2;
razn_h_mem[3628] = 132;
razn_h_mem[3629] = 8;
razn_h_mem[3630] = 138;
razn_h_mem[3631] = 14;
razn_h_mem[3632] = 144;
razn_h_mem[3633] = 20;
razn_h_mem[3634] = 150;
razn_h_mem[3635] = 26;
razn_h_mem[3636] = 156;
razn_h_mem[3637] = 32;
razn_h_mem[3638] = 162;
razn_h_mem[3639] = 38;
razn_h_mem[3640] = 168;
razn_h_mem[3641] = 44;
razn_h_mem[3642] = 174;
razn_h_mem[3643] = 50;
razn_h_mem[3644] = 180;
razn_h_mem[3645] = 56;
razn_h_mem[3646] = 186;
razn_h_mem[3647] = 62;
razn_h_mem[3648] = 192;
razn_h_mem[3649] = 68;
razn_h_mem[3650] = 198;
razn_h_mem[3651] = 74;
razn_h_mem[3652] = 204;
razn_h_mem[3653] = 80;
razn_h_mem[3654] = 210;
razn_h_mem[3655] = 86;
razn_h_mem[3656] = 216;
razn_h_mem[3657] = 92;
razn_h_mem[3658] = 222;
razn_h_mem[3659] = 98;
razn_h_mem[3660] = 228;
razn_h_mem[3661] = 104;
razn_h_mem[3662] = 234;
razn_h_mem[3663] = 110;
razn_h_mem[3664] = 240;
razn_h_mem[3665] = 116;
razn_h_mem[3666] = 246;
razn_h_mem[3667] = 122;
razn_h_mem[3668] = 252;
razn_h_mem[3669] = 128;
razn_h_mem[3670] = 4;
razn_h_mem[3671] = 134;
razn_h_mem[3672] = 10;
razn_h_mem[3673] = 140;
razn_h_mem[3674] = 16;
razn_h_mem[3675] = 146;
razn_h_mem[3676] = 22;
razn_h_mem[3677] = 152;
razn_h_mem[3678] = 28;
razn_h_mem[3679] = 158;
razn_h_mem[3680] = 34;
razn_h_mem[3681] = 164;
razn_h_mem[3682] = 40;
razn_h_mem[3683] = 170;
razn_h_mem[3684] = 46;
razn_h_mem[3685] = 176;
razn_h_mem[3686] = 52;
razn_h_mem[3687] = 182;
razn_h_mem[3688] = 58;
razn_h_mem[3689] = 188;
razn_h_mem[3690] = 64;
razn_h_mem[3691] = 194;
razn_h_mem[3692] = 70;
razn_h_mem[3693] = 200;
razn_h_mem[3694] = 76;
razn_h_mem[3695] = 206;
razn_h_mem[3696] = 82;
razn_h_mem[3697] = 212;
razn_h_mem[3698] = 88;
razn_h_mem[3699] = 218;
razn_h_mem[3700] = 94;
razn_h_mem[3701] = 224;
razn_h_mem[3702] = 100;
razn_h_mem[3703] = 230;
razn_h_mem[3704] = 106;
razn_h_mem[3705] = 236;
razn_h_mem[3706] = 112;
razn_h_mem[3707] = 242;
razn_h_mem[3708] = 118;
razn_h_mem[3709] = 248;
razn_h_mem[3710] = 124;
razn_h_mem[3711] = 255;
razn_h_mem[3712] = 0;
razn_h_mem[3713] = 130;
razn_h_mem[3714] = 6;
razn_h_mem[3715] = 136;
razn_h_mem[3716] = 12;
razn_h_mem[3717] = 142;
razn_h_mem[3718] = 18;
razn_h_mem[3719] = 148;
razn_h_mem[3720] = 24;
razn_h_mem[3721] = 154;
razn_h_mem[3722] = 30;
razn_h_mem[3723] = 160;
razn_h_mem[3724] = 36;
razn_h_mem[3725] = 166;
razn_h_mem[3726] = 42;
razn_h_mem[3727] = 172;
razn_h_mem[3728] = 48;
razn_h_mem[3729] = 178;
razn_h_mem[3730] = 54;
razn_h_mem[3731] = 184;
razn_h_mem[3732] = 60;
razn_h_mem[3733] = 190;
razn_h_mem[3734] = 66;
razn_h_mem[3735] = 196;
razn_h_mem[3736] = 72;
razn_h_mem[3737] = 202;
razn_h_mem[3738] = 78;
razn_h_mem[3739] = 208;
razn_h_mem[3740] = 84;
razn_h_mem[3741] = 214;
razn_h_mem[3742] = 90;
razn_h_mem[3743] = 220;
razn_h_mem[3744] = 96;
razn_h_mem[3745] = 226;
razn_h_mem[3746] = 102;
razn_h_mem[3747] = 232;
razn_h_mem[3748] = 108;
razn_h_mem[3749] = 238;
razn_h_mem[3750] = 114;
razn_h_mem[3751] = 244;
razn_h_mem[3752] = 120;
razn_h_mem[3753] = 250;
razn_h_mem[3754] = 126;
razn_h_mem[3755] = 2;
razn_h_mem[3756] = 132;
razn_h_mem[3757] = 8;
razn_h_mem[3758] = 138;
razn_h_mem[3759] = 14;
razn_h_mem[3760] = 144;
razn_h_mem[3761] = 20;
razn_h_mem[3762] = 150;
razn_h_mem[3763] = 26;
razn_h_mem[3764] = 156;
razn_h_mem[3765] = 32;
razn_h_mem[3766] = 162;
razn_h_mem[3767] = 38;
razn_h_mem[3768] = 168;
razn_h_mem[3769] = 44;
razn_h_mem[3770] = 174;
razn_h_mem[3771] = 50;
razn_h_mem[3772] = 180;
razn_h_mem[3773] = 56;
razn_h_mem[3774] = 186;
razn_h_mem[3775] = 62;
razn_h_mem[3776] = 192;
razn_h_mem[3777] = 68;
razn_h_mem[3778] = 198;
razn_h_mem[3779] = 74;
razn_h_mem[3780] = 204;
razn_h_mem[3781] = 80;
razn_h_mem[3782] = 210;
razn_h_mem[3783] = 86;
razn_h_mem[3784] = 216;
razn_h_mem[3785] = 92;
razn_h_mem[3786] = 222;
razn_h_mem[3787] = 98;
razn_h_mem[3788] = 228;
razn_h_mem[3789] = 104;
razn_h_mem[3790] = 234;
razn_h_mem[3791] = 110;
razn_h_mem[3792] = 240;
razn_h_mem[3793] = 116;
razn_h_mem[3794] = 246;
razn_h_mem[3795] = 122;
razn_h_mem[3796] = 252;
razn_h_mem[3797] = 128;
razn_h_mem[3798] = 4;
razn_h_mem[3799] = 134;
razn_h_mem[3800] = 10;
razn_h_mem[3801] = 140;
razn_h_mem[3802] = 16;
razn_h_mem[3803] = 146;
razn_h_mem[3804] = 22;
razn_h_mem[3805] = 152;
razn_h_mem[3806] = 28;
razn_h_mem[3807] = 158;
razn_h_mem[3808] = 34;
razn_h_mem[3809] = 164;
razn_h_mem[3810] = 40;
razn_h_mem[3811] = 170;
razn_h_mem[3812] = 46;
razn_h_mem[3813] = 176;
razn_h_mem[3814] = 52;
razn_h_mem[3815] = 182;
razn_h_mem[3816] = 58;
razn_h_mem[3817] = 188;
razn_h_mem[3818] = 64;
razn_h_mem[3819] = 194;
razn_h_mem[3820] = 70;
razn_h_mem[3821] = 200;
razn_h_mem[3822] = 76;
razn_h_mem[3823] = 206;
razn_h_mem[3824] = 82;
razn_h_mem[3825] = 212;
razn_h_mem[3826] = 88;
razn_h_mem[3827] = 218;
razn_h_mem[3828] = 94;
razn_h_mem[3829] = 224;
razn_h_mem[3830] = 100;
razn_h_mem[3831] = 230;
razn_h_mem[3832] = 106;
razn_h_mem[3833] = 236;
razn_h_mem[3834] = 112;
razn_h_mem[3835] = 242;
razn_h_mem[3836] = 118;
razn_h_mem[3837] = 248;
razn_h_mem[3838] = 124;
razn_h_mem[3839] = 255;
razn_h_mem[3840] = 0;
razn_h_mem[3841] = 130;
razn_h_mem[3842] = 6;
razn_h_mem[3843] = 136;
razn_h_mem[3844] = 12;
razn_h_mem[3845] = 142;
razn_h_mem[3846] = 18;
razn_h_mem[3847] = 148;
razn_h_mem[3848] = 24;
razn_h_mem[3849] = 154;
razn_h_mem[3850] = 30;
razn_h_mem[3851] = 160;
razn_h_mem[3852] = 36;
razn_h_mem[3853] = 166;
razn_h_mem[3854] = 42;
razn_h_mem[3855] = 172;
razn_h_mem[3856] = 48;
razn_h_mem[3857] = 178;
razn_h_mem[3858] = 54;
razn_h_mem[3859] = 184;
razn_h_mem[3860] = 60;
razn_h_mem[3861] = 190;
razn_h_mem[3862] = 66;
razn_h_mem[3863] = 196;
razn_h_mem[3864] = 72;
razn_h_mem[3865] = 202;
razn_h_mem[3866] = 78;
razn_h_mem[3867] = 208;
razn_h_mem[3868] = 84;
razn_h_mem[3869] = 214;
razn_h_mem[3870] = 90;
razn_h_mem[3871] = 220;
razn_h_mem[3872] = 96;
razn_h_mem[3873] = 226;
razn_h_mem[3874] = 102;
razn_h_mem[3875] = 232;
razn_h_mem[3876] = 108;
razn_h_mem[3877] = 238;
razn_h_mem[3878] = 114;
razn_h_mem[3879] = 244;
razn_h_mem[3880] = 120;
razn_h_mem[3881] = 250;
razn_h_mem[3882] = 126;
razn_h_mem[3883] = 2;
razn_h_mem[3884] = 132;
razn_h_mem[3885] = 8;
razn_h_mem[3886] = 138;
razn_h_mem[3887] = 14;
razn_h_mem[3888] = 144;
razn_h_mem[3889] = 20;
razn_h_mem[3890] = 150;
razn_h_mem[3891] = 26;
razn_h_mem[3892] = 156;
razn_h_mem[3893] = 32;
razn_h_mem[3894] = 162;
razn_h_mem[3895] = 38;
razn_h_mem[3896] = 168;
razn_h_mem[3897] = 44;
razn_h_mem[3898] = 174;
razn_h_mem[3899] = 50;
razn_h_mem[3900] = 180;
razn_h_mem[3901] = 56;
razn_h_mem[3902] = 186;
razn_h_mem[3903] = 62;
razn_h_mem[3904] = 192;
razn_h_mem[3905] = 68;
razn_h_mem[3906] = 198;
razn_h_mem[3907] = 74;
razn_h_mem[3908] = 204;
razn_h_mem[3909] = 80;
razn_h_mem[3910] = 210;
razn_h_mem[3911] = 86;
razn_h_mem[3912] = 216;
razn_h_mem[3913] = 92;
razn_h_mem[3914] = 222;
razn_h_mem[3915] = 98;
razn_h_mem[3916] = 228;
razn_h_mem[3917] = 104;
razn_h_mem[3918] = 234;
razn_h_mem[3919] = 110;
razn_h_mem[3920] = 240;
razn_h_mem[3921] = 116;
razn_h_mem[3922] = 246;
razn_h_mem[3923] = 122;
razn_h_mem[3924] = 252;
razn_h_mem[3925] = 128;
razn_h_mem[3926] = 4;
razn_h_mem[3927] = 134;
razn_h_mem[3928] = 10;
razn_h_mem[3929] = 140;
razn_h_mem[3930] = 16;
razn_h_mem[3931] = 146;
razn_h_mem[3932] = 22;
razn_h_mem[3933] = 152;
razn_h_mem[3934] = 28;
razn_h_mem[3935] = 158;
razn_h_mem[3936] = 34;
razn_h_mem[3937] = 164;
razn_h_mem[3938] = 40;
razn_h_mem[3939] = 170;
razn_h_mem[3940] = 46;
razn_h_mem[3941] = 176;
razn_h_mem[3942] = 52;
razn_h_mem[3943] = 182;
razn_h_mem[3944] = 58;
razn_h_mem[3945] = 188;
razn_h_mem[3946] = 64;
razn_h_mem[3947] = 194;
razn_h_mem[3948] = 70;
razn_h_mem[3949] = 200;
razn_h_mem[3950] = 76;
razn_h_mem[3951] = 206;
razn_h_mem[3952] = 82;
razn_h_mem[3953] = 212;
razn_h_mem[3954] = 88;
razn_h_mem[3955] = 218;
razn_h_mem[3956] = 94;
razn_h_mem[3957] = 224;
razn_h_mem[3958] = 100;
razn_h_mem[3959] = 230;
razn_h_mem[3960] = 106;
razn_h_mem[3961] = 236;
razn_h_mem[3962] = 112;
razn_h_mem[3963] = 242;
razn_h_mem[3964] = 118;
razn_h_mem[3965] = 248;
razn_h_mem[3966] = 124;
razn_h_mem[3967] = 255;
razn_h_mem[3968] = 0;
razn_h_mem[3969] = 130;
razn_h_mem[3970] = 6;
razn_h_mem[3971] = 136;
razn_h_mem[3972] = 12;
razn_h_mem[3973] = 142;
razn_h_mem[3974] = 18;
razn_h_mem[3975] = 148;
razn_h_mem[3976] = 24;
razn_h_mem[3977] = 154;
razn_h_mem[3978] = 30;
razn_h_mem[3979] = 160;
razn_h_mem[3980] = 36;
razn_h_mem[3981] = 166;
razn_h_mem[3982] = 42;
razn_h_mem[3983] = 172;
razn_h_mem[3984] = 48;
razn_h_mem[3985] = 178;
razn_h_mem[3986] = 54;
razn_h_mem[3987] = 184;
razn_h_mem[3988] = 60;
razn_h_mem[3989] = 190;
razn_h_mem[3990] = 66;
razn_h_mem[3991] = 196;
razn_h_mem[3992] = 72;
razn_h_mem[3993] = 202;
razn_h_mem[3994] = 78;
razn_h_mem[3995] = 208;
razn_h_mem[3996] = 84;
razn_h_mem[3997] = 214;
razn_h_mem[3998] = 90;
razn_h_mem[3999] = 220;
razn_h_mem[4000] = 96;
razn_h_mem[4001] = 226;
razn_h_mem[4002] = 102;
razn_h_mem[4003] = 232;
razn_h_mem[4004] = 108;
razn_h_mem[4005] = 238;
razn_h_mem[4006] = 114;
razn_h_mem[4007] = 244;
razn_h_mem[4008] = 120;
razn_h_mem[4009] = 250;
razn_h_mem[4010] = 126;
razn_h_mem[4011] = 2;
razn_h_mem[4012] = 132;
razn_h_mem[4013] = 8;
razn_h_mem[4014] = 138;
razn_h_mem[4015] = 14;
razn_h_mem[4016] = 144;
razn_h_mem[4017] = 20;
razn_h_mem[4018] = 150;
razn_h_mem[4019] = 26;
razn_h_mem[4020] = 156;
razn_h_mem[4021] = 32;
razn_h_mem[4022] = 162;
razn_h_mem[4023] = 38;
razn_h_mem[4024] = 168;
razn_h_mem[4025] = 44;
razn_h_mem[4026] = 174;
razn_h_mem[4027] = 50;
razn_h_mem[4028] = 180;
razn_h_mem[4029] = 56;
razn_h_mem[4030] = 186;
razn_h_mem[4031] = 62;
razn_h_mem[4032] = 192;
razn_h_mem[4033] = 68;
razn_h_mem[4034] = 198;
razn_h_mem[4035] = 74;
razn_h_mem[4036] = 204;
razn_h_mem[4037] = 80;
razn_h_mem[4038] = 210;
razn_h_mem[4039] = 86;
razn_h_mem[4040] = 216;
razn_h_mem[4041] = 92;
razn_h_mem[4042] = 222;
razn_h_mem[4043] = 98;
razn_h_mem[4044] = 228;
razn_h_mem[4045] = 104;
razn_h_mem[4046] = 234;
razn_h_mem[4047] = 110;
razn_h_mem[4048] = 240;
razn_h_mem[4049] = 116;
razn_h_mem[4050] = 246;
razn_h_mem[4051] = 122;
razn_h_mem[4052] = 252;
razn_h_mem[4053] = 128;
razn_h_mem[4054] = 4;
razn_h_mem[4055] = 134;
razn_h_mem[4056] = 10;
razn_h_mem[4057] = 140;
razn_h_mem[4058] = 16;
razn_h_mem[4059] = 146;
razn_h_mem[4060] = 22;
razn_h_mem[4061] = 152;
razn_h_mem[4062] = 28;
razn_h_mem[4063] = 158;
razn_h_mem[4064] = 34;
razn_h_mem[4065] = 164;
razn_h_mem[4066] = 40;
razn_h_mem[4067] = 170;
razn_h_mem[4068] = 46;
razn_h_mem[4069] = 176;
razn_h_mem[4070] = 52;
razn_h_mem[4071] = 182;
razn_h_mem[4072] = 58;
razn_h_mem[4073] = 188;
razn_h_mem[4074] = 64;
razn_h_mem[4075] = 194;
razn_h_mem[4076] = 70;
razn_h_mem[4077] = 200;
razn_h_mem[4078] = 76;
razn_h_mem[4079] = 206;
razn_h_mem[4080] = 82;
razn_h_mem[4081] = 212;
razn_h_mem[4082] = 88;
razn_h_mem[4083] = 218;
razn_h_mem[4084] = 94;
razn_h_mem[4085] = 224;
razn_h_mem[4086] = 100;
razn_h_mem[4087] = 230;
razn_h_mem[4088] = 106;
razn_h_mem[4089] = 236;
razn_h_mem[4090] = 112;
razn_h_mem[4091] = 242;
razn_h_mem[4092] = 118;
razn_h_mem[4093] = 248;
razn_h_mem[4094] = 124;
razn_h_mem[4095] = 255;
razn_h_mem[4096] = 0;
razn_h_mem[4097] = 130;
razn_h_mem[4098] = 6;
razn_h_mem[4099] = 136;
razn_h_mem[4100] = 12;
razn_h_mem[4101] = 142;
razn_h_mem[4102] = 18;
razn_h_mem[4103] = 148;
razn_h_mem[4104] = 24;
razn_h_mem[4105] = 154;
razn_h_mem[4106] = 30;
razn_h_mem[4107] = 160;
razn_h_mem[4108] = 36;
razn_h_mem[4109] = 166;
razn_h_mem[4110] = 42;
razn_h_mem[4111] = 172;
razn_h_mem[4112] = 48;
razn_h_mem[4113] = 178;
razn_h_mem[4114] = 54;
razn_h_mem[4115] = 184;
razn_h_mem[4116] = 60;
razn_h_mem[4117] = 190;
razn_h_mem[4118] = 66;
razn_h_mem[4119] = 196;
razn_h_mem[4120] = 72;
razn_h_mem[4121] = 202;
razn_h_mem[4122] = 78;
razn_h_mem[4123] = 208;
razn_h_mem[4124] = 84;
razn_h_mem[4125] = 214;
razn_h_mem[4126] = 90;
razn_h_mem[4127] = 220;
razn_h_mem[4128] = 96;
razn_h_mem[4129] = 226;
razn_h_mem[4130] = 102;
razn_h_mem[4131] = 232;
razn_h_mem[4132] = 108;
razn_h_mem[4133] = 238;
razn_h_mem[4134] = 114;
razn_h_mem[4135] = 244;
razn_h_mem[4136] = 120;
razn_h_mem[4137] = 250;
razn_h_mem[4138] = 126;
razn_h_mem[4139] = 2;
razn_h_mem[4140] = 132;
razn_h_mem[4141] = 8;
razn_h_mem[4142] = 138;
razn_h_mem[4143] = 14;
razn_h_mem[4144] = 144;
razn_h_mem[4145] = 20;
razn_h_mem[4146] = 150;
razn_h_mem[4147] = 26;
razn_h_mem[4148] = 156;
razn_h_mem[4149] = 32;
razn_h_mem[4150] = 162;
razn_h_mem[4151] = 38;
razn_h_mem[4152] = 168;
razn_h_mem[4153] = 44;
razn_h_mem[4154] = 174;
razn_h_mem[4155] = 50;
razn_h_mem[4156] = 180;
razn_h_mem[4157] = 56;
razn_h_mem[4158] = 186;
razn_h_mem[4159] = 62;
razn_h_mem[4160] = 192;
razn_h_mem[4161] = 68;
razn_h_mem[4162] = 198;
razn_h_mem[4163] = 74;
razn_h_mem[4164] = 204;
razn_h_mem[4165] = 80;
razn_h_mem[4166] = 210;
razn_h_mem[4167] = 86;
razn_h_mem[4168] = 216;
razn_h_mem[4169] = 92;
razn_h_mem[4170] = 222;
razn_h_mem[4171] = 98;
razn_h_mem[4172] = 228;
razn_h_mem[4173] = 104;
razn_h_mem[4174] = 234;
razn_h_mem[4175] = 110;
razn_h_mem[4176] = 240;
razn_h_mem[4177] = 116;
razn_h_mem[4178] = 246;
razn_h_mem[4179] = 122;
razn_h_mem[4180] = 252;
razn_h_mem[4181] = 128;
razn_h_mem[4182] = 4;
razn_h_mem[4183] = 134;
razn_h_mem[4184] = 10;
razn_h_mem[4185] = 140;
razn_h_mem[4186] = 16;
razn_h_mem[4187] = 146;
razn_h_mem[4188] = 22;
razn_h_mem[4189] = 152;
razn_h_mem[4190] = 28;
razn_h_mem[4191] = 158;
razn_h_mem[4192] = 34;
razn_h_mem[4193] = 164;
razn_h_mem[4194] = 40;
razn_h_mem[4195] = 170;
razn_h_mem[4196] = 46;
razn_h_mem[4197] = 176;
razn_h_mem[4198] = 52;
razn_h_mem[4199] = 182;
razn_h_mem[4200] = 58;
razn_h_mem[4201] = 188;
razn_h_mem[4202] = 64;
razn_h_mem[4203] = 194;
razn_h_mem[4204] = 70;
razn_h_mem[4205] = 200;
razn_h_mem[4206] = 76;
razn_h_mem[4207] = 206;
razn_h_mem[4208] = 82;
razn_h_mem[4209] = 212;
razn_h_mem[4210] = 88;
razn_h_mem[4211] = 218;
razn_h_mem[4212] = 94;
razn_h_mem[4213] = 224;
razn_h_mem[4214] = 100;
razn_h_mem[4215] = 230;
razn_h_mem[4216] = 106;
razn_h_mem[4217] = 236;
razn_h_mem[4218] = 112;
razn_h_mem[4219] = 242;
razn_h_mem[4220] = 118;
razn_h_mem[4221] = 248;
razn_h_mem[4222] = 124;
razn_h_mem[4223] = 255;
razn_h_mem[4224] = 0;
razn_h_mem[4225] = 130;
razn_h_mem[4226] = 6;
razn_h_mem[4227] = 136;
razn_h_mem[4228] = 12;
razn_h_mem[4229] = 142;
razn_h_mem[4230] = 18;
razn_h_mem[4231] = 148;
razn_h_mem[4232] = 24;
razn_h_mem[4233] = 154;
razn_h_mem[4234] = 30;
razn_h_mem[4235] = 160;
razn_h_mem[4236] = 36;
razn_h_mem[4237] = 166;
razn_h_mem[4238] = 42;
razn_h_mem[4239] = 172;
razn_h_mem[4240] = 48;
razn_h_mem[4241] = 178;
razn_h_mem[4242] = 54;
razn_h_mem[4243] = 184;
razn_h_mem[4244] = 60;
razn_h_mem[4245] = 190;
razn_h_mem[4246] = 66;
razn_h_mem[4247] = 196;
razn_h_mem[4248] = 72;
razn_h_mem[4249] = 202;
razn_h_mem[4250] = 78;
razn_h_mem[4251] = 208;
razn_h_mem[4252] = 84;
razn_h_mem[4253] = 214;
razn_h_mem[4254] = 90;
razn_h_mem[4255] = 220;
razn_h_mem[4256] = 96;
razn_h_mem[4257] = 226;
razn_h_mem[4258] = 102;
razn_h_mem[4259] = 232;
razn_h_mem[4260] = 108;
razn_h_mem[4261] = 238;
razn_h_mem[4262] = 114;
razn_h_mem[4263] = 244;
razn_h_mem[4264] = 120;
razn_h_mem[4265] = 250;
razn_h_mem[4266] = 126;
razn_h_mem[4267] = 2;
razn_h_mem[4268] = 132;
razn_h_mem[4269] = 8;
razn_h_mem[4270] = 138;
razn_h_mem[4271] = 14;
razn_h_mem[4272] = 144;
razn_h_mem[4273] = 20;
razn_h_mem[4274] = 150;
razn_h_mem[4275] = 26;
razn_h_mem[4276] = 156;
razn_h_mem[4277] = 32;
razn_h_mem[4278] = 162;
razn_h_mem[4279] = 38;
razn_h_mem[4280] = 168;
razn_h_mem[4281] = 44;
razn_h_mem[4282] = 174;
razn_h_mem[4283] = 50;
razn_h_mem[4284] = 180;
razn_h_mem[4285] = 56;
razn_h_mem[4286] = 186;
razn_h_mem[4287] = 62;
razn_h_mem[4288] = 192;
razn_h_mem[4289] = 68;
razn_h_mem[4290] = 198;
razn_h_mem[4291] = 74;
razn_h_mem[4292] = 204;
razn_h_mem[4293] = 80;
razn_h_mem[4294] = 210;
razn_h_mem[4295] = 86;
razn_h_mem[4296] = 216;
razn_h_mem[4297] = 92;
razn_h_mem[4298] = 222;
razn_h_mem[4299] = 98;
razn_h_mem[4300] = 228;
razn_h_mem[4301] = 104;
razn_h_mem[4302] = 234;
razn_h_mem[4303] = 110;
razn_h_mem[4304] = 240;
razn_h_mem[4305] = 116;
razn_h_mem[4306] = 246;
razn_h_mem[4307] = 122;
razn_h_mem[4308] = 252;
razn_h_mem[4309] = 128;
razn_h_mem[4310] = 4;
razn_h_mem[4311] = 134;
razn_h_mem[4312] = 10;
razn_h_mem[4313] = 140;
razn_h_mem[4314] = 16;
razn_h_mem[4315] = 146;
razn_h_mem[4316] = 22;
razn_h_mem[4317] = 152;
razn_h_mem[4318] = 28;
razn_h_mem[4319] = 158;
razn_h_mem[4320] = 34;
razn_h_mem[4321] = 164;
razn_h_mem[4322] = 40;
razn_h_mem[4323] = 170;
razn_h_mem[4324] = 46;
razn_h_mem[4325] = 176;
razn_h_mem[4326] = 52;
razn_h_mem[4327] = 182;
razn_h_mem[4328] = 58;
razn_h_mem[4329] = 188;
razn_h_mem[4330] = 64;
razn_h_mem[4331] = 194;
razn_h_mem[4332] = 70;
razn_h_mem[4333] = 200;
razn_h_mem[4334] = 76;
razn_h_mem[4335] = 206;
razn_h_mem[4336] = 82;
razn_h_mem[4337] = 212;
razn_h_mem[4338] = 88;
razn_h_mem[4339] = 218;
razn_h_mem[4340] = 94;
razn_h_mem[4341] = 224;
razn_h_mem[4342] = 100;
razn_h_mem[4343] = 230;
razn_h_mem[4344] = 106;
razn_h_mem[4345] = 236;
razn_h_mem[4346] = 112;
razn_h_mem[4347] = 242;
razn_h_mem[4348] = 118;
razn_h_mem[4349] = 248;
razn_h_mem[4350] = 124;
razn_h_mem[4351] = 255;
razn_h_mem[4352] = 0;
razn_h_mem[4353] = 130;
razn_h_mem[4354] = 6;
razn_h_mem[4355] = 136;
razn_h_mem[4356] = 12;
razn_h_mem[4357] = 142;
razn_h_mem[4358] = 18;
razn_h_mem[4359] = 148;
razn_h_mem[4360] = 24;
razn_h_mem[4361] = 154;
razn_h_mem[4362] = 30;
razn_h_mem[4363] = 160;
razn_h_mem[4364] = 36;
razn_h_mem[4365] = 166;
razn_h_mem[4366] = 42;
razn_h_mem[4367] = 172;
razn_h_mem[4368] = 48;
razn_h_mem[4369] = 178;
razn_h_mem[4370] = 54;
razn_h_mem[4371] = 184;
razn_h_mem[4372] = 60;
razn_h_mem[4373] = 190;
razn_h_mem[4374] = 66;
razn_h_mem[4375] = 196;
razn_h_mem[4376] = 72;
razn_h_mem[4377] = 202;
razn_h_mem[4378] = 78;
razn_h_mem[4379] = 208;
razn_h_mem[4380] = 84;
razn_h_mem[4381] = 214;
razn_h_mem[4382] = 90;
razn_h_mem[4383] = 220;
razn_h_mem[4384] = 96;
razn_h_mem[4385] = 226;
razn_h_mem[4386] = 102;
razn_h_mem[4387] = 232;
razn_h_mem[4388] = 108;
razn_h_mem[4389] = 238;
razn_h_mem[4390] = 114;
razn_h_mem[4391] = 244;
razn_h_mem[4392] = 120;
razn_h_mem[4393] = 250;
razn_h_mem[4394] = 126;
razn_h_mem[4395] = 2;
razn_h_mem[4396] = 132;
razn_h_mem[4397] = 8;
razn_h_mem[4398] = 138;
razn_h_mem[4399] = 14;
razn_h_mem[4400] = 144;
razn_h_mem[4401] = 20;
razn_h_mem[4402] = 150;
razn_h_mem[4403] = 26;
razn_h_mem[4404] = 156;
razn_h_mem[4405] = 32;
razn_h_mem[4406] = 162;
razn_h_mem[4407] = 38;
razn_h_mem[4408] = 168;
razn_h_mem[4409] = 44;
razn_h_mem[4410] = 174;
razn_h_mem[4411] = 50;
razn_h_mem[4412] = 180;
razn_h_mem[4413] = 56;
razn_h_mem[4414] = 186;
razn_h_mem[4415] = 62;
razn_h_mem[4416] = 192;
razn_h_mem[4417] = 68;
razn_h_mem[4418] = 198;
razn_h_mem[4419] = 74;
razn_h_mem[4420] = 204;
razn_h_mem[4421] = 80;
razn_h_mem[4422] = 210;
razn_h_mem[4423] = 86;
razn_h_mem[4424] = 216;
razn_h_mem[4425] = 92;
razn_h_mem[4426] = 222;
razn_h_mem[4427] = 98;
razn_h_mem[4428] = 228;
razn_h_mem[4429] = 104;
razn_h_mem[4430] = 234;
razn_h_mem[4431] = 110;
razn_h_mem[4432] = 240;
razn_h_mem[4433] = 116;
razn_h_mem[4434] = 246;
razn_h_mem[4435] = 122;
razn_h_mem[4436] = 252;
razn_h_mem[4437] = 128;
razn_h_mem[4438] = 4;
razn_h_mem[4439] = 134;
razn_h_mem[4440] = 10;
razn_h_mem[4441] = 140;
razn_h_mem[4442] = 16;
razn_h_mem[4443] = 146;
razn_h_mem[4444] = 22;
razn_h_mem[4445] = 152;
razn_h_mem[4446] = 28;
razn_h_mem[4447] = 158;
razn_h_mem[4448] = 34;
razn_h_mem[4449] = 164;
razn_h_mem[4450] = 40;
razn_h_mem[4451] = 170;
razn_h_mem[4452] = 46;
razn_h_mem[4453] = 176;
razn_h_mem[4454] = 52;
razn_h_mem[4455] = 182;
razn_h_mem[4456] = 58;
razn_h_mem[4457] = 188;
razn_h_mem[4458] = 64;
razn_h_mem[4459] = 194;
razn_h_mem[4460] = 70;
razn_h_mem[4461] = 200;
razn_h_mem[4462] = 76;
razn_h_mem[4463] = 206;
razn_h_mem[4464] = 82;
razn_h_mem[4465] = 212;
razn_h_mem[4466] = 88;
razn_h_mem[4467] = 218;
razn_h_mem[4468] = 94;
razn_h_mem[4469] = 224;
razn_h_mem[4470] = 100;
razn_h_mem[4471] = 230;
razn_h_mem[4472] = 106;
razn_h_mem[4473] = 236;
razn_h_mem[4474] = 112;
razn_h_mem[4475] = 242;
razn_h_mem[4476] = 118;
razn_h_mem[4477] = 248;
razn_h_mem[4478] = 124;
razn_h_mem[4479] = 255;
razn_h_mem[4480] = 0;
razn_h_mem[4481] = 130;
razn_h_mem[4482] = 6;
razn_h_mem[4483] = 136;
razn_h_mem[4484] = 12;
razn_h_mem[4485] = 142;
razn_h_mem[4486] = 18;
razn_h_mem[4487] = 148;
razn_h_mem[4488] = 24;
razn_h_mem[4489] = 154;
razn_h_mem[4490] = 30;
razn_h_mem[4491] = 160;
razn_h_mem[4492] = 36;
razn_h_mem[4493] = 166;
razn_h_mem[4494] = 42;
razn_h_mem[4495] = 172;
razn_h_mem[4496] = 48;
razn_h_mem[4497] = 178;
razn_h_mem[4498] = 54;
razn_h_mem[4499] = 184;
razn_h_mem[4500] = 60;
razn_h_mem[4501] = 190;
razn_h_mem[4502] = 66;
razn_h_mem[4503] = 196;
razn_h_mem[4504] = 72;
razn_h_mem[4505] = 202;
razn_h_mem[4506] = 78;
razn_h_mem[4507] = 208;
razn_h_mem[4508] = 84;
razn_h_mem[4509] = 214;
razn_h_mem[4510] = 90;
razn_h_mem[4511] = 220;
razn_h_mem[4512] = 96;
razn_h_mem[4513] = 226;
razn_h_mem[4514] = 102;
razn_h_mem[4515] = 232;
razn_h_mem[4516] = 108;
razn_h_mem[4517] = 238;
razn_h_mem[4518] = 114;
razn_h_mem[4519] = 244;
razn_h_mem[4520] = 120;
razn_h_mem[4521] = 250;
razn_h_mem[4522] = 126;
razn_h_mem[4523] = 2;
razn_h_mem[4524] = 132;
razn_h_mem[4525] = 8;
razn_h_mem[4526] = 138;
razn_h_mem[4527] = 14;
razn_h_mem[4528] = 144;
razn_h_mem[4529] = 20;
razn_h_mem[4530] = 150;
razn_h_mem[4531] = 26;
razn_h_mem[4532] = 156;
razn_h_mem[4533] = 32;
razn_h_mem[4534] = 162;
razn_h_mem[4535] = 38;
razn_h_mem[4536] = 168;
razn_h_mem[4537] = 44;
razn_h_mem[4538] = 174;
razn_h_mem[4539] = 50;
razn_h_mem[4540] = 180;
razn_h_mem[4541] = 56;
razn_h_mem[4542] = 186;
razn_h_mem[4543] = 62;
razn_h_mem[4544] = 192;
razn_h_mem[4545] = 68;
razn_h_mem[4546] = 198;
razn_h_mem[4547] = 74;
razn_h_mem[4548] = 204;
razn_h_mem[4549] = 80;
razn_h_mem[4550] = 210;
razn_h_mem[4551] = 86;
razn_h_mem[4552] = 216;
razn_h_mem[4553] = 92;
razn_h_mem[4554] = 222;
razn_h_mem[4555] = 98;
razn_h_mem[4556] = 228;
razn_h_mem[4557] = 104;
razn_h_mem[4558] = 234;
razn_h_mem[4559] = 110;
razn_h_mem[4560] = 240;
razn_h_mem[4561] = 116;
razn_h_mem[4562] = 246;
razn_h_mem[4563] = 122;
razn_h_mem[4564] = 252;
razn_h_mem[4565] = 128;
razn_h_mem[4566] = 4;
razn_h_mem[4567] = 134;
razn_h_mem[4568] = 10;
razn_h_mem[4569] = 140;
razn_h_mem[4570] = 16;
razn_h_mem[4571] = 146;
razn_h_mem[4572] = 22;
razn_h_mem[4573] = 152;
razn_h_mem[4574] = 28;
razn_h_mem[4575] = 158;
razn_h_mem[4576] = 34;
razn_h_mem[4577] = 164;
razn_h_mem[4578] = 40;
razn_h_mem[4579] = 170;
razn_h_mem[4580] = 46;
razn_h_mem[4581] = 176;
razn_h_mem[4582] = 52;
razn_h_mem[4583] = 182;
razn_h_mem[4584] = 58;
razn_h_mem[4585] = 188;
razn_h_mem[4586] = 64;
razn_h_mem[4587] = 194;
razn_h_mem[4588] = 70;
razn_h_mem[4589] = 200;
razn_h_mem[4590] = 76;
razn_h_mem[4591] = 206;
razn_h_mem[4592] = 82;
razn_h_mem[4593] = 212;
razn_h_mem[4594] = 88;
razn_h_mem[4595] = 218;
razn_h_mem[4596] = 94;
razn_h_mem[4597] = 224;
razn_h_mem[4598] = 100;
razn_h_mem[4599] = 230;
razn_h_mem[4600] = 106;
razn_h_mem[4601] = 236;
razn_h_mem[4602] = 112;
razn_h_mem[4603] = 242;
razn_h_mem[4604] = 118;
razn_h_mem[4605] = 248;
razn_h_mem[4606] = 124;
razn_h_mem[4607] = 255;
razn_h_mem[4608] = 0;
razn_h_mem[4609] = 130;
razn_h_mem[4610] = 6;
razn_h_mem[4611] = 136;
razn_h_mem[4612] = 12;
razn_h_mem[4613] = 142;
razn_h_mem[4614] = 18;
razn_h_mem[4615] = 148;
razn_h_mem[4616] = 24;
razn_h_mem[4617] = 154;
razn_h_mem[4618] = 30;
razn_h_mem[4619] = 160;
razn_h_mem[4620] = 36;
razn_h_mem[4621] = 166;
razn_h_mem[4622] = 42;
razn_h_mem[4623] = 172;
razn_h_mem[4624] = 48;
razn_h_mem[4625] = 178;
razn_h_mem[4626] = 54;
razn_h_mem[4627] = 184;
razn_h_mem[4628] = 60;
razn_h_mem[4629] = 190;
razn_h_mem[4630] = 66;
razn_h_mem[4631] = 196;
razn_h_mem[4632] = 72;
razn_h_mem[4633] = 202;
razn_h_mem[4634] = 78;
razn_h_mem[4635] = 208;
razn_h_mem[4636] = 84;
razn_h_mem[4637] = 214;
razn_h_mem[4638] = 90;
razn_h_mem[4639] = 220;
razn_h_mem[4640] = 96;
razn_h_mem[4641] = 226;
razn_h_mem[4642] = 102;
razn_h_mem[4643] = 232;
razn_h_mem[4644] = 108;
razn_h_mem[4645] = 238;
razn_h_mem[4646] = 114;
razn_h_mem[4647] = 244;
razn_h_mem[4648] = 120;
razn_h_mem[4649] = 250;
razn_h_mem[4650] = 126;
razn_h_mem[4651] = 2;
razn_h_mem[4652] = 132;
razn_h_mem[4653] = 8;
razn_h_mem[4654] = 138;
razn_h_mem[4655] = 14;
razn_h_mem[4656] = 144;
razn_h_mem[4657] = 20;
razn_h_mem[4658] = 150;
razn_h_mem[4659] = 26;
razn_h_mem[4660] = 156;
razn_h_mem[4661] = 32;
razn_h_mem[4662] = 162;
razn_h_mem[4663] = 38;
razn_h_mem[4664] = 168;
razn_h_mem[4665] = 44;
razn_h_mem[4666] = 174;
razn_h_mem[4667] = 50;
razn_h_mem[4668] = 180;
razn_h_mem[4669] = 56;
razn_h_mem[4670] = 186;
razn_h_mem[4671] = 62;
razn_h_mem[4672] = 192;
razn_h_mem[4673] = 68;
razn_h_mem[4674] = 198;
razn_h_mem[4675] = 74;
razn_h_mem[4676] = 204;
razn_h_mem[4677] = 80;
razn_h_mem[4678] = 210;
razn_h_mem[4679] = 86;
razn_h_mem[4680] = 216;
razn_h_mem[4681] = 92;
razn_h_mem[4682] = 222;
razn_h_mem[4683] = 98;
razn_h_mem[4684] = 228;
razn_h_mem[4685] = 104;
razn_h_mem[4686] = 234;
razn_h_mem[4687] = 110;
razn_h_mem[4688] = 240;
razn_h_mem[4689] = 116;
razn_h_mem[4690] = 246;
razn_h_mem[4691] = 122;
razn_h_mem[4692] = 252;
razn_h_mem[4693] = 128;
razn_h_mem[4694] = 4;
razn_h_mem[4695] = 134;
razn_h_mem[4696] = 10;
razn_h_mem[4697] = 140;
razn_h_mem[4698] = 16;
razn_h_mem[4699] = 146;
razn_h_mem[4700] = 22;
razn_h_mem[4701] = 152;
razn_h_mem[4702] = 28;
razn_h_mem[4703] = 158;
razn_h_mem[4704] = 34;
razn_h_mem[4705] = 164;
razn_h_mem[4706] = 40;
razn_h_mem[4707] = 170;
razn_h_mem[4708] = 46;
razn_h_mem[4709] = 176;
razn_h_mem[4710] = 52;
razn_h_mem[4711] = 182;
razn_h_mem[4712] = 58;
razn_h_mem[4713] = 188;
razn_h_mem[4714] = 64;
razn_h_mem[4715] = 194;
razn_h_mem[4716] = 70;
razn_h_mem[4717] = 200;
razn_h_mem[4718] = 76;
razn_h_mem[4719] = 206;
razn_h_mem[4720] = 82;
razn_h_mem[4721] = 212;
razn_h_mem[4722] = 88;
razn_h_mem[4723] = 218;
razn_h_mem[4724] = 94;
razn_h_mem[4725] = 224;
razn_h_mem[4726] = 100;
razn_h_mem[4727] = 230;
razn_h_mem[4728] = 106;
razn_h_mem[4729] = 236;
razn_h_mem[4730] = 112;
razn_h_mem[4731] = 242;
razn_h_mem[4732] = 118;
razn_h_mem[4733] = 248;
razn_h_mem[4734] = 124;
razn_h_mem[4735] = 255;
razn_h_mem[4736] = 0;
razn_h_mem[4737] = 130;
razn_h_mem[4738] = 6;
razn_h_mem[4739] = 136;
razn_h_mem[4740] = 12;
razn_h_mem[4741] = 142;
razn_h_mem[4742] = 18;
razn_h_mem[4743] = 148;
razn_h_mem[4744] = 24;
razn_h_mem[4745] = 154;
razn_h_mem[4746] = 30;
razn_h_mem[4747] = 160;
razn_h_mem[4748] = 36;
razn_h_mem[4749] = 166;
razn_h_mem[4750] = 42;
razn_h_mem[4751] = 172;
razn_h_mem[4752] = 48;
razn_h_mem[4753] = 178;
razn_h_mem[4754] = 54;
razn_h_mem[4755] = 184;
razn_h_mem[4756] = 60;
razn_h_mem[4757] = 190;
razn_h_mem[4758] = 66;
razn_h_mem[4759] = 196;
razn_h_mem[4760] = 72;
razn_h_mem[4761] = 202;
razn_h_mem[4762] = 78;
razn_h_mem[4763] = 208;
razn_h_mem[4764] = 84;
razn_h_mem[4765] = 214;
razn_h_mem[4766] = 90;
razn_h_mem[4767] = 220;
razn_h_mem[4768] = 96;
razn_h_mem[4769] = 226;
razn_h_mem[4770] = 102;
razn_h_mem[4771] = 232;
razn_h_mem[4772] = 108;
razn_h_mem[4773] = 238;
razn_h_mem[4774] = 114;
razn_h_mem[4775] = 244;
razn_h_mem[4776] = 120;
razn_h_mem[4777] = 250;
razn_h_mem[4778] = 126;
razn_h_mem[4779] = 2;
razn_h_mem[4780] = 132;
razn_h_mem[4781] = 8;
razn_h_mem[4782] = 138;
razn_h_mem[4783] = 14;
razn_h_mem[4784] = 144;
razn_h_mem[4785] = 20;
razn_h_mem[4786] = 150;
razn_h_mem[4787] = 26;
razn_h_mem[4788] = 156;
razn_h_mem[4789] = 32;
razn_h_mem[4790] = 162;
razn_h_mem[4791] = 38;
razn_h_mem[4792] = 168;
razn_h_mem[4793] = 44;
razn_h_mem[4794] = 174;
razn_h_mem[4795] = 50;
razn_h_mem[4796] = 180;
razn_h_mem[4797] = 56;
razn_h_mem[4798] = 186;
razn_h_mem[4799] = 62;
razn_h_mem[4800] = 192;
razn_h_mem[4801] = 68;
razn_h_mem[4802] = 198;
razn_h_mem[4803] = 74;
razn_h_mem[4804] = 204;
razn_h_mem[4805] = 80;
razn_h_mem[4806] = 210;
razn_h_mem[4807] = 86;
razn_h_mem[4808] = 216;
razn_h_mem[4809] = 92;
razn_h_mem[4810] = 222;
razn_h_mem[4811] = 98;
razn_h_mem[4812] = 228;
razn_h_mem[4813] = 104;
razn_h_mem[4814] = 234;
razn_h_mem[4815] = 110;
razn_h_mem[4816] = 240;
razn_h_mem[4817] = 116;
razn_h_mem[4818] = 246;
razn_h_mem[4819] = 122;
razn_h_mem[4820] = 252;
razn_h_mem[4821] = 128;
razn_h_mem[4822] = 4;
razn_h_mem[4823] = 134;
razn_h_mem[4824] = 10;
razn_h_mem[4825] = 140;
razn_h_mem[4826] = 16;
razn_h_mem[4827] = 146;
razn_h_mem[4828] = 22;
razn_h_mem[4829] = 152;
razn_h_mem[4830] = 28;
razn_h_mem[4831] = 158;
razn_h_mem[4832] = 34;
razn_h_mem[4833] = 164;
razn_h_mem[4834] = 40;
razn_h_mem[4835] = 170;
razn_h_mem[4836] = 46;
razn_h_mem[4837] = 176;
razn_h_mem[4838] = 52;
razn_h_mem[4839] = 182;
razn_h_mem[4840] = 58;
razn_h_mem[4841] = 188;
razn_h_mem[4842] = 64;
razn_h_mem[4843] = 194;
razn_h_mem[4844] = 70;
razn_h_mem[4845] = 200;
razn_h_mem[4846] = 76;
razn_h_mem[4847] = 206;
razn_h_mem[4848] = 82;
razn_h_mem[4849] = 212;
razn_h_mem[4850] = 88;
razn_h_mem[4851] = 218;
razn_h_mem[4852] = 94;
razn_h_mem[4853] = 224;
razn_h_mem[4854] = 100;
razn_h_mem[4855] = 230;
razn_h_mem[4856] = 106;
razn_h_mem[4857] = 236;
razn_h_mem[4858] = 112;
razn_h_mem[4859] = 242;
razn_h_mem[4860] = 118;
razn_h_mem[4861] = 248;
razn_h_mem[4862] = 124;
razn_h_mem[4863] = 255;
razn_h_mem[4864] = 0;
razn_h_mem[4865] = 130;
razn_h_mem[4866] = 6;
razn_h_mem[4867] = 136;
razn_h_mem[4868] = 12;
razn_h_mem[4869] = 142;
razn_h_mem[4870] = 18;
razn_h_mem[4871] = 148;
razn_h_mem[4872] = 24;
razn_h_mem[4873] = 154;
razn_h_mem[4874] = 30;
razn_h_mem[4875] = 160;
razn_h_mem[4876] = 36;
razn_h_mem[4877] = 166;
razn_h_mem[4878] = 42;
razn_h_mem[4879] = 172;
razn_h_mem[4880] = 48;
razn_h_mem[4881] = 178;
razn_h_mem[4882] = 54;
razn_h_mem[4883] = 184;
razn_h_mem[4884] = 60;
razn_h_mem[4885] = 190;
razn_h_mem[4886] = 66;
razn_h_mem[4887] = 196;
razn_h_mem[4888] = 72;
razn_h_mem[4889] = 202;
razn_h_mem[4890] = 78;
razn_h_mem[4891] = 208;
razn_h_mem[4892] = 84;
razn_h_mem[4893] = 214;
razn_h_mem[4894] = 90;
razn_h_mem[4895] = 220;
razn_h_mem[4896] = 96;
razn_h_mem[4897] = 226;
razn_h_mem[4898] = 102;
razn_h_mem[4899] = 232;
razn_h_mem[4900] = 108;
razn_h_mem[4901] = 238;
razn_h_mem[4902] = 114;
razn_h_mem[4903] = 244;
razn_h_mem[4904] = 120;
razn_h_mem[4905] = 250;
razn_h_mem[4906] = 126;
razn_h_mem[4907] = 2;
razn_h_mem[4908] = 132;
razn_h_mem[4909] = 8;
razn_h_mem[4910] = 138;
razn_h_mem[4911] = 14;
razn_h_mem[4912] = 144;
razn_h_mem[4913] = 20;
razn_h_mem[4914] = 150;
razn_h_mem[4915] = 26;
razn_h_mem[4916] = 156;
razn_h_mem[4917] = 32;
razn_h_mem[4918] = 162;
razn_h_mem[4919] = 38;
razn_h_mem[4920] = 168;
razn_h_mem[4921] = 44;
razn_h_mem[4922] = 174;
razn_h_mem[4923] = 50;
razn_h_mem[4924] = 180;
razn_h_mem[4925] = 56;
razn_h_mem[4926] = 186;
razn_h_mem[4927] = 62;
razn_h_mem[4928] = 192;
razn_h_mem[4929] = 68;
razn_h_mem[4930] = 198;
razn_h_mem[4931] = 74;
razn_h_mem[4932] = 204;
razn_h_mem[4933] = 80;
razn_h_mem[4934] = 210;
razn_h_mem[4935] = 86;
razn_h_mem[4936] = 216;
razn_h_mem[4937] = 92;
razn_h_mem[4938] = 222;
razn_h_mem[4939] = 98;
razn_h_mem[4940] = 228;
razn_h_mem[4941] = 104;
razn_h_mem[4942] = 234;
razn_h_mem[4943] = 110;
razn_h_mem[4944] = 240;
razn_h_mem[4945] = 116;
razn_h_mem[4946] = 246;
razn_h_mem[4947] = 122;
razn_h_mem[4948] = 252;
razn_h_mem[4949] = 128;
razn_h_mem[4950] = 4;
razn_h_mem[4951] = 134;
razn_h_mem[4952] = 10;
razn_h_mem[4953] = 140;
razn_h_mem[4954] = 16;
razn_h_mem[4955] = 146;
razn_h_mem[4956] = 22;
razn_h_mem[4957] = 152;
razn_h_mem[4958] = 28;
razn_h_mem[4959] = 158;
razn_h_mem[4960] = 34;
razn_h_mem[4961] = 164;
razn_h_mem[4962] = 40;
razn_h_mem[4963] = 170;
razn_h_mem[4964] = 46;
razn_h_mem[4965] = 176;
razn_h_mem[4966] = 52;
razn_h_mem[4967] = 182;
razn_h_mem[4968] = 58;
razn_h_mem[4969] = 188;
razn_h_mem[4970] = 64;
razn_h_mem[4971] = 194;
razn_h_mem[4972] = 70;
razn_h_mem[4973] = 200;
razn_h_mem[4974] = 76;
razn_h_mem[4975] = 206;
razn_h_mem[4976] = 82;
razn_h_mem[4977] = 212;
razn_h_mem[4978] = 88;
razn_h_mem[4979] = 218;
razn_h_mem[4980] = 94;
razn_h_mem[4981] = 224;
razn_h_mem[4982] = 100;
razn_h_mem[4983] = 230;
razn_h_mem[4984] = 106;
razn_h_mem[4985] = 236;
razn_h_mem[4986] = 112;
razn_h_mem[4987] = 242;
razn_h_mem[4988] = 118;
razn_h_mem[4989] = 248;
razn_h_mem[4990] = 124;
razn_h_mem[4991] = 255;
razn_h_mem[4992] = 0;
razn_h_mem[4993] = 130;
razn_h_mem[4994] = 6;
razn_h_mem[4995] = 136;
razn_h_mem[4996] = 12;
razn_h_mem[4997] = 142;
razn_h_mem[4998] = 18;
razn_h_mem[4999] = 148;
razn_h_mem[5000] = 24;
razn_h_mem[5001] = 154;
razn_h_mem[5002] = 30;
razn_h_mem[5003] = 160;
razn_h_mem[5004] = 36;
razn_h_mem[5005] = 166;
razn_h_mem[5006] = 42;
razn_h_mem[5007] = 172;
razn_h_mem[5008] = 48;
razn_h_mem[5009] = 178;
razn_h_mem[5010] = 54;
razn_h_mem[5011] = 184;
razn_h_mem[5012] = 60;
razn_h_mem[5013] = 190;
razn_h_mem[5014] = 66;
razn_h_mem[5015] = 196;
razn_h_mem[5016] = 72;
razn_h_mem[5017] = 202;
razn_h_mem[5018] = 78;
razn_h_mem[5019] = 208;
razn_h_mem[5020] = 84;
razn_h_mem[5021] = 214;
razn_h_mem[5022] = 90;
razn_h_mem[5023] = 220;
razn_h_mem[5024] = 96;
razn_h_mem[5025] = 226;
razn_h_mem[5026] = 102;
razn_h_mem[5027] = 232;
razn_h_mem[5028] = 108;
razn_h_mem[5029] = 238;
razn_h_mem[5030] = 114;
razn_h_mem[5031] = 244;
razn_h_mem[5032] = 120;
razn_h_mem[5033] = 250;
razn_h_mem[5034] = 126;
razn_h_mem[5035] = 2;
razn_h_mem[5036] = 132;
razn_h_mem[5037] = 8;
razn_h_mem[5038] = 138;
razn_h_mem[5039] = 14;
razn_h_mem[5040] = 144;
razn_h_mem[5041] = 20;
razn_h_mem[5042] = 150;
razn_h_mem[5043] = 26;
razn_h_mem[5044] = 156;
razn_h_mem[5045] = 32;
razn_h_mem[5046] = 162;
razn_h_mem[5047] = 38;
razn_h_mem[5048] = 168;
razn_h_mem[5049] = 44;
razn_h_mem[5050] = 174;
razn_h_mem[5051] = 50;
razn_h_mem[5052] = 180;
razn_h_mem[5053] = 56;
razn_h_mem[5054] = 186;
razn_h_mem[5055] = 62;
razn_h_mem[5056] = 192;
razn_h_mem[5057] = 68;
razn_h_mem[5058] = 198;
razn_h_mem[5059] = 74;
razn_h_mem[5060] = 204;
razn_h_mem[5061] = 80;
razn_h_mem[5062] = 210;
razn_h_mem[5063] = 86;
razn_h_mem[5064] = 216;
razn_h_mem[5065] = 92;
razn_h_mem[5066] = 222;
razn_h_mem[5067] = 98;
razn_h_mem[5068] = 228;
razn_h_mem[5069] = 104;
razn_h_mem[5070] = 234;
razn_h_mem[5071] = 110;
razn_h_mem[5072] = 240;
razn_h_mem[5073] = 116;
razn_h_mem[5074] = 246;
razn_h_mem[5075] = 122;
razn_h_mem[5076] = 252;
razn_h_mem[5077] = 128;
razn_h_mem[5078] = 4;
razn_h_mem[5079] = 134;
razn_h_mem[5080] = 10;
razn_h_mem[5081] = 140;
razn_h_mem[5082] = 16;
razn_h_mem[5083] = 146;
razn_h_mem[5084] = 22;
razn_h_mem[5085] = 152;
razn_h_mem[5086] = 28;
razn_h_mem[5087] = 158;
razn_h_mem[5088] = 34;
razn_h_mem[5089] = 164;
razn_h_mem[5090] = 40;
razn_h_mem[5091] = 170;
razn_h_mem[5092] = 46;
razn_h_mem[5093] = 176;
razn_h_mem[5094] = 52;
razn_h_mem[5095] = 182;
razn_h_mem[5096] = 58;
razn_h_mem[5097] = 188;
razn_h_mem[5098] = 64;
razn_h_mem[5099] = 194;
razn_h_mem[5100] = 70;
razn_h_mem[5101] = 200;
razn_h_mem[5102] = 76;
razn_h_mem[5103] = 206;
razn_h_mem[5104] = 82;
razn_h_mem[5105] = 212;
razn_h_mem[5106] = 88;
razn_h_mem[5107] = 218;
razn_h_mem[5108] = 94;
razn_h_mem[5109] = 224;
razn_h_mem[5110] = 100;
razn_h_mem[5111] = 230;
razn_h_mem[5112] = 106;
razn_h_mem[5113] = 236;
razn_h_mem[5114] = 112;
razn_h_mem[5115] = 242;
razn_h_mem[5116] = 118;
razn_h_mem[5117] = 248;
razn_h_mem[5118] = 124;
razn_h_mem[5119] = 255;
razn_h_mem[5120] = 0;
razn_h_mem[5121] = 130;
razn_h_mem[5122] = 6;
razn_h_mem[5123] = 136;
razn_h_mem[5124] = 12;
razn_h_mem[5125] = 142;
razn_h_mem[5126] = 18;
razn_h_mem[5127] = 148;
razn_h_mem[5128] = 24;
razn_h_mem[5129] = 154;
razn_h_mem[5130] = 30;
razn_h_mem[5131] = 160;
razn_h_mem[5132] = 36;
razn_h_mem[5133] = 166;
razn_h_mem[5134] = 42;
razn_h_mem[5135] = 172;
razn_h_mem[5136] = 48;
razn_h_mem[5137] = 178;
razn_h_mem[5138] = 54;
razn_h_mem[5139] = 184;
razn_h_mem[5140] = 60;
razn_h_mem[5141] = 190;
razn_h_mem[5142] = 66;
razn_h_mem[5143] = 196;
razn_h_mem[5144] = 72;
razn_h_mem[5145] = 202;
razn_h_mem[5146] = 78;
razn_h_mem[5147] = 208;
razn_h_mem[5148] = 84;
razn_h_mem[5149] = 214;
razn_h_mem[5150] = 90;
razn_h_mem[5151] = 220;
razn_h_mem[5152] = 96;
razn_h_mem[5153] = 226;
razn_h_mem[5154] = 102;
razn_h_mem[5155] = 232;
razn_h_mem[5156] = 108;
razn_h_mem[5157] = 238;
razn_h_mem[5158] = 114;
razn_h_mem[5159] = 244;
razn_h_mem[5160] = 120;
razn_h_mem[5161] = 250;
razn_h_mem[5162] = 126;
razn_h_mem[5163] = 2;
razn_h_mem[5164] = 132;
razn_h_mem[5165] = 8;
razn_h_mem[5166] = 138;
razn_h_mem[5167] = 14;
razn_h_mem[5168] = 144;
razn_h_mem[5169] = 20;
razn_h_mem[5170] = 150;
razn_h_mem[5171] = 26;
razn_h_mem[5172] = 156;
razn_h_mem[5173] = 32;
razn_h_mem[5174] = 162;
razn_h_mem[5175] = 38;
razn_h_mem[5176] = 168;
razn_h_mem[5177] = 44;
razn_h_mem[5178] = 174;
razn_h_mem[5179] = 50;
razn_h_mem[5180] = 180;
razn_h_mem[5181] = 56;
razn_h_mem[5182] = 186;
razn_h_mem[5183] = 62;
razn_h_mem[5184] = 192;
razn_h_mem[5185] = 68;
razn_h_mem[5186] = 198;
razn_h_mem[5187] = 74;
razn_h_mem[5188] = 204;
razn_h_mem[5189] = 80;
razn_h_mem[5190] = 210;
razn_h_mem[5191] = 86;
razn_h_mem[5192] = 216;
razn_h_mem[5193] = 92;
razn_h_mem[5194] = 222;
razn_h_mem[5195] = 98;
razn_h_mem[5196] = 228;
razn_h_mem[5197] = 104;
razn_h_mem[5198] = 234;
razn_h_mem[5199] = 110;
razn_h_mem[5200] = 240;
razn_h_mem[5201] = 116;
razn_h_mem[5202] = 246;
razn_h_mem[5203] = 122;
razn_h_mem[5204] = 252;
razn_h_mem[5205] = 128;
razn_h_mem[5206] = 4;
razn_h_mem[5207] = 134;
razn_h_mem[5208] = 10;
razn_h_mem[5209] = 140;
razn_h_mem[5210] = 16;
razn_h_mem[5211] = 146;
razn_h_mem[5212] = 22;
razn_h_mem[5213] = 152;
razn_h_mem[5214] = 28;
razn_h_mem[5215] = 158;
razn_h_mem[5216] = 34;
razn_h_mem[5217] = 164;
razn_h_mem[5218] = 40;
razn_h_mem[5219] = 170;
razn_h_mem[5220] = 46;
razn_h_mem[5221] = 176;
razn_h_mem[5222] = 52;
razn_h_mem[5223] = 182;
razn_h_mem[5224] = 58;
razn_h_mem[5225] = 188;
razn_h_mem[5226] = 64;
razn_h_mem[5227] = 194;
razn_h_mem[5228] = 70;
razn_h_mem[5229] = 200;
razn_h_mem[5230] = 76;
razn_h_mem[5231] = 206;
razn_h_mem[5232] = 82;
razn_h_mem[5233] = 212;
razn_h_mem[5234] = 88;
razn_h_mem[5235] = 218;
razn_h_mem[5236] = 94;
razn_h_mem[5237] = 224;
razn_h_mem[5238] = 100;
razn_h_mem[5239] = 230;
razn_h_mem[5240] = 106;
razn_h_mem[5241] = 236;
razn_h_mem[5242] = 112;
razn_h_mem[5243] = 242;
razn_h_mem[5244] = 118;
razn_h_mem[5245] = 248;
razn_h_mem[5246] = 124;
razn_h_mem[5247] = 255;
razn_h_mem[5248] = 0;
razn_h_mem[5249] = 130;
razn_h_mem[5250] = 6;
razn_h_mem[5251] = 136;
razn_h_mem[5252] = 12;
razn_h_mem[5253] = 142;
razn_h_mem[5254] = 18;
razn_h_mem[5255] = 148;
razn_h_mem[5256] = 24;
razn_h_mem[5257] = 154;
razn_h_mem[5258] = 30;
razn_h_mem[5259] = 160;
razn_h_mem[5260] = 36;
razn_h_mem[5261] = 166;
razn_h_mem[5262] = 42;
razn_h_mem[5263] = 172;
razn_h_mem[5264] = 48;
razn_h_mem[5265] = 178;
razn_h_mem[5266] = 54;
razn_h_mem[5267] = 184;
razn_h_mem[5268] = 60;
razn_h_mem[5269] = 190;
razn_h_mem[5270] = 66;
razn_h_mem[5271] = 196;
razn_h_mem[5272] = 72;
razn_h_mem[5273] = 202;
razn_h_mem[5274] = 78;
razn_h_mem[5275] = 208;
razn_h_mem[5276] = 84;
razn_h_mem[5277] = 214;
razn_h_mem[5278] = 90;
razn_h_mem[5279] = 220;
razn_h_mem[5280] = 96;
razn_h_mem[5281] = 226;
razn_h_mem[5282] = 102;
razn_h_mem[5283] = 232;
razn_h_mem[5284] = 108;
razn_h_mem[5285] = 238;
razn_h_mem[5286] = 114;
razn_h_mem[5287] = 244;
razn_h_mem[5288] = 120;
razn_h_mem[5289] = 250;
razn_h_mem[5290] = 126;
razn_h_mem[5291] = 2;
razn_h_mem[5292] = 132;
razn_h_mem[5293] = 8;
razn_h_mem[5294] = 138;
razn_h_mem[5295] = 14;
razn_h_mem[5296] = 144;
razn_h_mem[5297] = 20;
razn_h_mem[5298] = 150;
razn_h_mem[5299] = 26;
razn_h_mem[5300] = 156;
razn_h_mem[5301] = 32;
razn_h_mem[5302] = 162;
razn_h_mem[5303] = 38;
razn_h_mem[5304] = 168;
razn_h_mem[5305] = 44;
razn_h_mem[5306] = 174;
razn_h_mem[5307] = 50;
razn_h_mem[5308] = 180;
razn_h_mem[5309] = 56;
razn_h_mem[5310] = 186;
razn_h_mem[5311] = 62;
razn_h_mem[5312] = 192;
razn_h_mem[5313] = 68;
razn_h_mem[5314] = 198;
razn_h_mem[5315] = 74;
razn_h_mem[5316] = 204;
razn_h_mem[5317] = 80;
razn_h_mem[5318] = 210;
razn_h_mem[5319] = 86;
razn_h_mem[5320] = 216;
razn_h_mem[5321] = 92;
razn_h_mem[5322] = 222;
razn_h_mem[5323] = 98;
razn_h_mem[5324] = 228;
razn_h_mem[5325] = 104;
razn_h_mem[5326] = 234;
razn_h_mem[5327] = 110;
razn_h_mem[5328] = 240;
razn_h_mem[5329] = 116;
razn_h_mem[5330] = 246;
razn_h_mem[5331] = 122;
razn_h_mem[5332] = 252;
razn_h_mem[5333] = 128;
razn_h_mem[5334] = 4;
razn_h_mem[5335] = 134;
razn_h_mem[5336] = 10;
razn_h_mem[5337] = 140;
razn_h_mem[5338] = 16;
razn_h_mem[5339] = 146;
razn_h_mem[5340] = 22;
razn_h_mem[5341] = 152;
razn_h_mem[5342] = 28;
razn_h_mem[5343] = 158;
razn_h_mem[5344] = 34;
razn_h_mem[5345] = 164;
razn_h_mem[5346] = 40;
razn_h_mem[5347] = 170;
razn_h_mem[5348] = 46;
razn_h_mem[5349] = 176;
razn_h_mem[5350] = 52;
razn_h_mem[5351] = 182;
razn_h_mem[5352] = 58;
razn_h_mem[5353] = 188;
razn_h_mem[5354] = 64;
razn_h_mem[5355] = 194;
razn_h_mem[5356] = 70;
razn_h_mem[5357] = 200;
razn_h_mem[5358] = 76;
razn_h_mem[5359] = 206;
razn_h_mem[5360] = 82;
razn_h_mem[5361] = 212;
razn_h_mem[5362] = 88;
razn_h_mem[5363] = 218;
razn_h_mem[5364] = 94;
razn_h_mem[5365] = 224;
razn_h_mem[5366] = 100;
razn_h_mem[5367] = 230;
razn_h_mem[5368] = 106;
razn_h_mem[5369] = 236;
razn_h_mem[5370] = 112;
razn_h_mem[5371] = 242;
razn_h_mem[5372] = 118;
razn_h_mem[5373] = 248;
razn_h_mem[5374] = 124;
razn_h_mem[5375] = 255;
razn_h_mem[5376] = 0;
razn_h_mem[5377] = 130;
razn_h_mem[5378] = 6;
razn_h_mem[5379] = 136;
razn_h_mem[5380] = 12;
razn_h_mem[5381] = 142;
razn_h_mem[5382] = 18;
razn_h_mem[5383] = 148;
razn_h_mem[5384] = 24;
razn_h_mem[5385] = 154;
razn_h_mem[5386] = 30;
razn_h_mem[5387] = 160;
razn_h_mem[5388] = 36;
razn_h_mem[5389] = 166;
razn_h_mem[5390] = 42;
razn_h_mem[5391] = 172;
razn_h_mem[5392] = 48;
razn_h_mem[5393] = 178;
razn_h_mem[5394] = 54;
razn_h_mem[5395] = 184;
razn_h_mem[5396] = 60;
razn_h_mem[5397] = 190;
razn_h_mem[5398] = 66;
razn_h_mem[5399] = 196;
razn_h_mem[5400] = 72;
razn_h_mem[5401] = 202;
razn_h_mem[5402] = 78;
razn_h_mem[5403] = 208;
razn_h_mem[5404] = 84;
razn_h_mem[5405] = 214;
razn_h_mem[5406] = 90;
razn_h_mem[5407] = 220;
razn_h_mem[5408] = 96;
razn_h_mem[5409] = 226;
razn_h_mem[5410] = 102;
razn_h_mem[5411] = 232;
razn_h_mem[5412] = 108;
razn_h_mem[5413] = 238;
razn_h_mem[5414] = 114;
razn_h_mem[5415] = 244;
razn_h_mem[5416] = 120;
razn_h_mem[5417] = 250;
razn_h_mem[5418] = 126;
razn_h_mem[5419] = 2;
razn_h_mem[5420] = 132;
razn_h_mem[5421] = 8;
razn_h_mem[5422] = 138;
razn_h_mem[5423] = 14;
razn_h_mem[5424] = 144;
razn_h_mem[5425] = 20;
razn_h_mem[5426] = 150;
razn_h_mem[5427] = 26;
razn_h_mem[5428] = 156;
razn_h_mem[5429] = 32;
razn_h_mem[5430] = 162;
razn_h_mem[5431] = 38;
razn_h_mem[5432] = 168;
razn_h_mem[5433] = 44;
razn_h_mem[5434] = 174;
razn_h_mem[5435] = 50;
razn_h_mem[5436] = 180;
razn_h_mem[5437] = 56;
razn_h_mem[5438] = 186;
razn_h_mem[5439] = 62;
razn_h_mem[5440] = 192;
razn_h_mem[5441] = 68;
razn_h_mem[5442] = 198;
razn_h_mem[5443] = 74;
razn_h_mem[5444] = 204;
razn_h_mem[5445] = 80;
razn_h_mem[5446] = 210;
razn_h_mem[5447] = 86;
razn_h_mem[5448] = 216;
razn_h_mem[5449] = 92;
razn_h_mem[5450] = 222;
razn_h_mem[5451] = 98;
razn_h_mem[5452] = 228;
razn_h_mem[5453] = 104;
razn_h_mem[5454] = 234;
razn_h_mem[5455] = 110;
razn_h_mem[5456] = 240;
razn_h_mem[5457] = 116;
razn_h_mem[5458] = 246;
razn_h_mem[5459] = 122;
razn_h_mem[5460] = 252;
razn_h_mem[5461] = 128;
razn_h_mem[5462] = 4;
razn_h_mem[5463] = 134;
razn_h_mem[5464] = 10;
razn_h_mem[5465] = 140;
razn_h_mem[5466] = 16;
razn_h_mem[5467] = 146;
razn_h_mem[5468] = 22;
razn_h_mem[5469] = 152;
razn_h_mem[5470] = 28;
razn_h_mem[5471] = 158;
razn_h_mem[5472] = 34;
razn_h_mem[5473] = 164;
razn_h_mem[5474] = 40;
razn_h_mem[5475] = 170;
razn_h_mem[5476] = 46;
razn_h_mem[5477] = 176;
razn_h_mem[5478] = 52;
razn_h_mem[5479] = 182;
razn_h_mem[5480] = 58;
razn_h_mem[5481] = 188;
razn_h_mem[5482] = 64;
razn_h_mem[5483] = 194;
razn_h_mem[5484] = 70;
razn_h_mem[5485] = 200;
razn_h_mem[5486] = 76;
razn_h_mem[5487] = 206;
razn_h_mem[5488] = 82;
razn_h_mem[5489] = 212;
razn_h_mem[5490] = 88;
razn_h_mem[5491] = 218;
razn_h_mem[5492] = 94;
razn_h_mem[5493] = 224;
razn_h_mem[5494] = 100;
razn_h_mem[5495] = 230;
razn_h_mem[5496] = 106;
razn_h_mem[5497] = 236;
razn_h_mem[5498] = 112;
razn_h_mem[5499] = 242;
razn_h_mem[5500] = 118;
razn_h_mem[5501] = 248;
razn_h_mem[5502] = 124;
razn_h_mem[5503] = 255;
razn_h_mem[5504] = 0;
razn_h_mem[5505] = 130;
razn_h_mem[5506] = 6;
razn_h_mem[5507] = 136;
razn_h_mem[5508] = 12;
razn_h_mem[5509] = 142;
razn_h_mem[5510] = 18;
razn_h_mem[5511] = 148;
razn_h_mem[5512] = 24;
razn_h_mem[5513] = 154;
razn_h_mem[5514] = 30;
razn_h_mem[5515] = 160;
razn_h_mem[5516] = 36;
razn_h_mem[5517] = 166;
razn_h_mem[5518] = 42;
razn_h_mem[5519] = 172;
razn_h_mem[5520] = 48;
razn_h_mem[5521] = 178;
razn_h_mem[5522] = 54;
razn_h_mem[5523] = 184;
razn_h_mem[5524] = 60;
razn_h_mem[5525] = 190;
razn_h_mem[5526] = 66;
razn_h_mem[5527] = 196;
razn_h_mem[5528] = 72;
razn_h_mem[5529] = 202;
razn_h_mem[5530] = 78;
razn_h_mem[5531] = 208;
razn_h_mem[5532] = 84;
razn_h_mem[5533] = 214;
razn_h_mem[5534] = 90;
razn_h_mem[5535] = 220;
razn_h_mem[5536] = 96;
razn_h_mem[5537] = 226;
razn_h_mem[5538] = 102;
razn_h_mem[5539] = 232;
razn_h_mem[5540] = 108;
razn_h_mem[5541] = 238;
razn_h_mem[5542] = 114;
razn_h_mem[5543] = 244;
razn_h_mem[5544] = 120;
razn_h_mem[5545] = 250;
razn_h_mem[5546] = 126;
razn_h_mem[5547] = 2;
razn_h_mem[5548] = 132;
razn_h_mem[5549] = 8;
razn_h_mem[5550] = 138;
razn_h_mem[5551] = 14;
razn_h_mem[5552] = 144;
razn_h_mem[5553] = 20;
razn_h_mem[5554] = 150;
razn_h_mem[5555] = 26;
razn_h_mem[5556] = 156;
razn_h_mem[5557] = 32;
razn_h_mem[5558] = 162;
razn_h_mem[5559] = 38;
razn_h_mem[5560] = 168;
razn_h_mem[5561] = 44;
razn_h_mem[5562] = 174;
razn_h_mem[5563] = 50;
razn_h_mem[5564] = 180;
razn_h_mem[5565] = 56;
razn_h_mem[5566] = 186;
razn_h_mem[5567] = 62;
razn_h_mem[5568] = 192;
razn_h_mem[5569] = 68;
razn_h_mem[5570] = 198;
razn_h_mem[5571] = 74;
razn_h_mem[5572] = 204;
razn_h_mem[5573] = 80;
razn_h_mem[5574] = 210;
razn_h_mem[5575] = 86;
razn_h_mem[5576] = 216;
razn_h_mem[5577] = 92;
razn_h_mem[5578] = 222;
razn_h_mem[5579] = 98;
razn_h_mem[5580] = 228;
razn_h_mem[5581] = 104;
razn_h_mem[5582] = 234;
razn_h_mem[5583] = 110;
razn_h_mem[5584] = 240;
razn_h_mem[5585] = 116;
razn_h_mem[5586] = 246;
razn_h_mem[5587] = 122;
razn_h_mem[5588] = 252;
razn_h_mem[5589] = 128;
razn_h_mem[5590] = 4;
razn_h_mem[5591] = 134;
razn_h_mem[5592] = 10;
razn_h_mem[5593] = 140;
razn_h_mem[5594] = 16;
razn_h_mem[5595] = 146;
razn_h_mem[5596] = 22;
razn_h_mem[5597] = 152;
razn_h_mem[5598] = 28;
razn_h_mem[5599] = 158;
razn_h_mem[5600] = 34;
razn_h_mem[5601] = 164;
razn_h_mem[5602] = 40;
razn_h_mem[5603] = 170;
razn_h_mem[5604] = 46;
razn_h_mem[5605] = 176;
razn_h_mem[5606] = 52;
razn_h_mem[5607] = 182;
razn_h_mem[5608] = 58;
razn_h_mem[5609] = 188;
razn_h_mem[5610] = 64;
razn_h_mem[5611] = 194;
razn_h_mem[5612] = 70;
razn_h_mem[5613] = 200;
razn_h_mem[5614] = 76;
razn_h_mem[5615] = 206;
razn_h_mem[5616] = 82;
razn_h_mem[5617] = 212;
razn_h_mem[5618] = 88;
razn_h_mem[5619] = 218;
razn_h_mem[5620] = 94;
razn_h_mem[5621] = 224;
razn_h_mem[5622] = 100;
razn_h_mem[5623] = 230;
razn_h_mem[5624] = 106;
razn_h_mem[5625] = 236;
razn_h_mem[5626] = 112;
razn_h_mem[5627] = 242;
razn_h_mem[5628] = 118;
razn_h_mem[5629] = 248;
razn_h_mem[5630] = 124;
razn_h_mem[5631] = 255;
razn_h_mem[5632] = 0;
razn_h_mem[5633] = 130;
razn_h_mem[5634] = 6;
razn_h_mem[5635] = 136;
razn_h_mem[5636] = 12;
razn_h_mem[5637] = 142;
razn_h_mem[5638] = 18;
razn_h_mem[5639] = 148;
razn_h_mem[5640] = 24;
razn_h_mem[5641] = 154;
razn_h_mem[5642] = 30;
razn_h_mem[5643] = 160;
razn_h_mem[5644] = 36;
razn_h_mem[5645] = 166;
razn_h_mem[5646] = 42;
razn_h_mem[5647] = 172;
razn_h_mem[5648] = 48;
razn_h_mem[5649] = 178;
razn_h_mem[5650] = 54;
razn_h_mem[5651] = 184;
razn_h_mem[5652] = 60;
razn_h_mem[5653] = 190;
razn_h_mem[5654] = 66;
razn_h_mem[5655] = 196;
razn_h_mem[5656] = 72;
razn_h_mem[5657] = 202;
razn_h_mem[5658] = 78;
razn_h_mem[5659] = 208;
razn_h_mem[5660] = 84;
razn_h_mem[5661] = 214;
razn_h_mem[5662] = 90;
razn_h_mem[5663] = 220;
razn_h_mem[5664] = 96;
razn_h_mem[5665] = 226;
razn_h_mem[5666] = 102;
razn_h_mem[5667] = 232;
razn_h_mem[5668] = 108;
razn_h_mem[5669] = 238;
razn_h_mem[5670] = 114;
razn_h_mem[5671] = 244;
razn_h_mem[5672] = 120;
razn_h_mem[5673] = 250;
razn_h_mem[5674] = 126;
razn_h_mem[5675] = 2;
razn_h_mem[5676] = 132;
razn_h_mem[5677] = 8;
razn_h_mem[5678] = 138;
razn_h_mem[5679] = 14;
razn_h_mem[5680] = 144;
razn_h_mem[5681] = 20;
razn_h_mem[5682] = 150;
razn_h_mem[5683] = 26;
razn_h_mem[5684] = 156;
razn_h_mem[5685] = 32;
razn_h_mem[5686] = 162;
razn_h_mem[5687] = 38;
razn_h_mem[5688] = 168;
razn_h_mem[5689] = 44;
razn_h_mem[5690] = 174;
razn_h_mem[5691] = 50;
razn_h_mem[5692] = 180;
razn_h_mem[5693] = 56;
razn_h_mem[5694] = 186;
razn_h_mem[5695] = 62;
razn_h_mem[5696] = 192;
razn_h_mem[5697] = 68;
razn_h_mem[5698] = 198;
razn_h_mem[5699] = 74;
razn_h_mem[5700] = 204;
razn_h_mem[5701] = 80;
razn_h_mem[5702] = 210;
razn_h_mem[5703] = 86;
razn_h_mem[5704] = 216;
razn_h_mem[5705] = 92;
razn_h_mem[5706] = 222;
razn_h_mem[5707] = 98;
razn_h_mem[5708] = 228;
razn_h_mem[5709] = 104;
razn_h_mem[5710] = 234;
razn_h_mem[5711] = 110;
razn_h_mem[5712] = 240;
razn_h_mem[5713] = 116;
razn_h_mem[5714] = 246;
razn_h_mem[5715] = 122;
razn_h_mem[5716] = 252;
razn_h_mem[5717] = 128;
razn_h_mem[5718] = 4;
razn_h_mem[5719] = 134;
razn_h_mem[5720] = 10;
razn_h_mem[5721] = 140;
razn_h_mem[5722] = 16;
razn_h_mem[5723] = 146;
razn_h_mem[5724] = 22;
razn_h_mem[5725] = 152;
razn_h_mem[5726] = 28;
razn_h_mem[5727] = 158;
razn_h_mem[5728] = 34;
razn_h_mem[5729] = 164;
razn_h_mem[5730] = 40;
razn_h_mem[5731] = 170;
razn_h_mem[5732] = 46;
razn_h_mem[5733] = 176;
razn_h_mem[5734] = 52;
razn_h_mem[5735] = 182;
razn_h_mem[5736] = 58;
razn_h_mem[5737] = 188;
razn_h_mem[5738] = 64;
razn_h_mem[5739] = 194;
razn_h_mem[5740] = 70;
razn_h_mem[5741] = 200;
razn_h_mem[5742] = 76;
razn_h_mem[5743] = 206;
razn_h_mem[5744] = 82;
razn_h_mem[5745] = 212;
razn_h_mem[5746] = 88;
razn_h_mem[5747] = 218;
razn_h_mem[5748] = 94;
razn_h_mem[5749] = 224;
razn_h_mem[5750] = 100;
razn_h_mem[5751] = 230;
razn_h_mem[5752] = 106;
razn_h_mem[5753] = 236;
razn_h_mem[5754] = 112;
razn_h_mem[5755] = 242;
razn_h_mem[5756] = 118;
razn_h_mem[5757] = 248;
razn_h_mem[5758] = 124;
razn_h_mem[5759] = 255;
razn_h_mem[5760] = 0;
razn_h_mem[5761] = 130;
razn_h_mem[5762] = 6;
razn_h_mem[5763] = 136;
razn_h_mem[5764] = 12;
razn_h_mem[5765] = 142;
razn_h_mem[5766] = 18;
razn_h_mem[5767] = 148;
razn_h_mem[5768] = 24;
razn_h_mem[5769] = 154;
razn_h_mem[5770] = 30;
razn_h_mem[5771] = 160;
razn_h_mem[5772] = 36;
razn_h_mem[5773] = 166;
razn_h_mem[5774] = 42;
razn_h_mem[5775] = 172;
razn_h_mem[5776] = 48;
razn_h_mem[5777] = 178;
razn_h_mem[5778] = 54;
razn_h_mem[5779] = 184;
razn_h_mem[5780] = 60;
razn_h_mem[5781] = 190;
razn_h_mem[5782] = 66;
razn_h_mem[5783] = 196;
razn_h_mem[5784] = 72;
razn_h_mem[5785] = 202;
razn_h_mem[5786] = 78;
razn_h_mem[5787] = 208;
razn_h_mem[5788] = 84;
razn_h_mem[5789] = 214;
razn_h_mem[5790] = 90;
razn_h_mem[5791] = 220;
razn_h_mem[5792] = 96;
razn_h_mem[5793] = 226;
razn_h_mem[5794] = 102;
razn_h_mem[5795] = 232;
razn_h_mem[5796] = 108;
razn_h_mem[5797] = 238;
razn_h_mem[5798] = 114;
razn_h_mem[5799] = 244;
razn_h_mem[5800] = 120;
razn_h_mem[5801] = 250;
razn_h_mem[5802] = 126;
razn_h_mem[5803] = 2;
razn_h_mem[5804] = 132;
razn_h_mem[5805] = 8;
razn_h_mem[5806] = 138;
razn_h_mem[5807] = 14;
razn_h_mem[5808] = 144;
razn_h_mem[5809] = 20;
razn_h_mem[5810] = 150;
razn_h_mem[5811] = 26;
razn_h_mem[5812] = 156;
razn_h_mem[5813] = 32;
razn_h_mem[5814] = 162;
razn_h_mem[5815] = 38;
razn_h_mem[5816] = 168;
razn_h_mem[5817] = 44;
razn_h_mem[5818] = 174;
razn_h_mem[5819] = 50;
razn_h_mem[5820] = 180;
razn_h_mem[5821] = 56;
razn_h_mem[5822] = 186;
razn_h_mem[5823] = 62;
razn_h_mem[5824] = 192;
razn_h_mem[5825] = 68;
razn_h_mem[5826] = 198;
razn_h_mem[5827] = 74;
razn_h_mem[5828] = 204;
razn_h_mem[5829] = 80;
razn_h_mem[5830] = 210;
razn_h_mem[5831] = 86;
razn_h_mem[5832] = 216;
razn_h_mem[5833] = 92;
razn_h_mem[5834] = 222;
razn_h_mem[5835] = 98;
razn_h_mem[5836] = 228;
razn_h_mem[5837] = 104;
razn_h_mem[5838] = 234;
razn_h_mem[5839] = 110;
razn_h_mem[5840] = 240;
razn_h_mem[5841] = 116;
razn_h_mem[5842] = 246;
razn_h_mem[5843] = 122;
razn_h_mem[5844] = 252;
razn_h_mem[5845] = 128;
razn_h_mem[5846] = 4;
razn_h_mem[5847] = 134;
razn_h_mem[5848] = 10;
razn_h_mem[5849] = 140;
razn_h_mem[5850] = 16;
razn_h_mem[5851] = 146;
razn_h_mem[5852] = 22;
razn_h_mem[5853] = 152;
razn_h_mem[5854] = 28;
razn_h_mem[5855] = 158;
razn_h_mem[5856] = 34;
razn_h_mem[5857] = 164;
razn_h_mem[5858] = 40;
razn_h_mem[5859] = 170;
razn_h_mem[5860] = 46;
razn_h_mem[5861] = 176;
razn_h_mem[5862] = 52;
razn_h_mem[5863] = 182;
razn_h_mem[5864] = 58;
razn_h_mem[5865] = 188;
razn_h_mem[5866] = 64;
razn_h_mem[5867] = 194;
razn_h_mem[5868] = 70;
razn_h_mem[5869] = 200;
razn_h_mem[5870] = 76;
razn_h_mem[5871] = 206;
razn_h_mem[5872] = 82;
razn_h_mem[5873] = 212;
razn_h_mem[5874] = 88;
razn_h_mem[5875] = 218;
razn_h_mem[5876] = 94;
razn_h_mem[5877] = 224;
razn_h_mem[5878] = 100;
razn_h_mem[5879] = 230;
razn_h_mem[5880] = 106;
razn_h_mem[5881] = 236;
razn_h_mem[5882] = 112;
razn_h_mem[5883] = 242;
razn_h_mem[5884] = 118;
razn_h_mem[5885] = 248;
razn_h_mem[5886] = 124;
razn_h_mem[5887] = 255;
razn_h_mem[5888] = 0;
razn_h_mem[5889] = 130;
razn_h_mem[5890] = 6;
razn_h_mem[5891] = 136;
razn_h_mem[5892] = 12;
razn_h_mem[5893] = 142;
razn_h_mem[5894] = 18;
razn_h_mem[5895] = 148;
razn_h_mem[5896] = 24;
razn_h_mem[5897] = 154;
razn_h_mem[5898] = 30;
razn_h_mem[5899] = 160;
razn_h_mem[5900] = 36;
razn_h_mem[5901] = 166;
razn_h_mem[5902] = 42;
razn_h_mem[5903] = 172;
razn_h_mem[5904] = 48;
razn_h_mem[5905] = 178;
razn_h_mem[5906] = 54;
razn_h_mem[5907] = 184;
razn_h_mem[5908] = 60;
razn_h_mem[5909] = 190;
razn_h_mem[5910] = 66;
razn_h_mem[5911] = 196;
razn_h_mem[5912] = 72;
razn_h_mem[5913] = 202;
razn_h_mem[5914] = 78;
razn_h_mem[5915] = 208;
razn_h_mem[5916] = 84;
razn_h_mem[5917] = 214;
razn_h_mem[5918] = 90;
razn_h_mem[5919] = 220;
razn_h_mem[5920] = 96;
razn_h_mem[5921] = 226;
razn_h_mem[5922] = 102;
razn_h_mem[5923] = 232;
razn_h_mem[5924] = 108;
razn_h_mem[5925] = 238;
razn_h_mem[5926] = 114;
razn_h_mem[5927] = 244;
razn_h_mem[5928] = 120;
razn_h_mem[5929] = 250;
razn_h_mem[5930] = 126;
razn_h_mem[5931] = 2;
razn_h_mem[5932] = 132;
razn_h_mem[5933] = 8;
razn_h_mem[5934] = 138;
razn_h_mem[5935] = 14;
razn_h_mem[5936] = 144;
razn_h_mem[5937] = 20;
razn_h_mem[5938] = 150;
razn_h_mem[5939] = 26;
razn_h_mem[5940] = 156;
razn_h_mem[5941] = 32;
razn_h_mem[5942] = 162;
razn_h_mem[5943] = 38;
razn_h_mem[5944] = 168;
razn_h_mem[5945] = 44;
razn_h_mem[5946] = 174;
razn_h_mem[5947] = 50;
razn_h_mem[5948] = 180;
razn_h_mem[5949] = 56;
razn_h_mem[5950] = 186;
razn_h_mem[5951] = 62;
razn_h_mem[5952] = 192;
razn_h_mem[5953] = 68;
razn_h_mem[5954] = 198;
razn_h_mem[5955] = 74;
razn_h_mem[5956] = 204;
razn_h_mem[5957] = 80;
razn_h_mem[5958] = 210;
razn_h_mem[5959] = 86;
razn_h_mem[5960] = 216;
razn_h_mem[5961] = 92;
razn_h_mem[5962] = 222;
razn_h_mem[5963] = 98;
razn_h_mem[5964] = 228;
razn_h_mem[5965] = 104;
razn_h_mem[5966] = 234;
razn_h_mem[5967] = 110;
razn_h_mem[5968] = 240;
razn_h_mem[5969] = 116;
razn_h_mem[5970] = 246;
razn_h_mem[5971] = 122;
razn_h_mem[5972] = 252;
razn_h_mem[5973] = 128;
razn_h_mem[5974] = 4;
razn_h_mem[5975] = 134;
razn_h_mem[5976] = 10;
razn_h_mem[5977] = 140;
razn_h_mem[5978] = 16;
razn_h_mem[5979] = 146;
razn_h_mem[5980] = 22;
razn_h_mem[5981] = 152;
razn_h_mem[5982] = 28;
razn_h_mem[5983] = 158;
razn_h_mem[5984] = 34;
razn_h_mem[5985] = 164;
razn_h_mem[5986] = 40;
razn_h_mem[5987] = 170;
razn_h_mem[5988] = 46;
razn_h_mem[5989] = 176;
razn_h_mem[5990] = 52;
razn_h_mem[5991] = 182;
razn_h_mem[5992] = 58;
razn_h_mem[5993] = 188;
razn_h_mem[5994] = 64;
razn_h_mem[5995] = 194;
razn_h_mem[5996] = 70;
razn_h_mem[5997] = 200;
razn_h_mem[5998] = 76;
razn_h_mem[5999] = 206;
razn_h_mem[6000] = 82;
razn_h_mem[6001] = 212;
razn_h_mem[6002] = 88;
razn_h_mem[6003] = 218;
razn_h_mem[6004] = 94;
razn_h_mem[6005] = 224;
razn_h_mem[6006] = 100;
razn_h_mem[6007] = 230;
razn_h_mem[6008] = 106;
razn_h_mem[6009] = 236;
razn_h_mem[6010] = 112;
razn_h_mem[6011] = 242;
razn_h_mem[6012] = 118;
razn_h_mem[6013] = 248;
razn_h_mem[6014] = 124;
razn_h_mem[6015] = 255;
razn_h_mem[6016] = 0;
razn_h_mem[6017] = 130;
razn_h_mem[6018] = 6;
razn_h_mem[6019] = 136;
razn_h_mem[6020] = 12;
razn_h_mem[6021] = 142;
razn_h_mem[6022] = 18;
razn_h_mem[6023] = 148;
razn_h_mem[6024] = 24;
razn_h_mem[6025] = 154;
razn_h_mem[6026] = 30;
razn_h_mem[6027] = 160;
razn_h_mem[6028] = 36;
razn_h_mem[6029] = 166;
razn_h_mem[6030] = 42;
razn_h_mem[6031] = 172;
razn_h_mem[6032] = 48;
razn_h_mem[6033] = 178;
razn_h_mem[6034] = 54;
razn_h_mem[6035] = 184;
razn_h_mem[6036] = 60;
razn_h_mem[6037] = 190;
razn_h_mem[6038] = 66;
razn_h_mem[6039] = 196;
razn_h_mem[6040] = 72;
razn_h_mem[6041] = 202;
razn_h_mem[6042] = 78;
razn_h_mem[6043] = 208;
razn_h_mem[6044] = 84;
razn_h_mem[6045] = 214;
razn_h_mem[6046] = 90;
razn_h_mem[6047] = 220;
razn_h_mem[6048] = 96;
razn_h_mem[6049] = 226;
razn_h_mem[6050] = 102;
razn_h_mem[6051] = 232;
razn_h_mem[6052] = 108;
razn_h_mem[6053] = 238;
razn_h_mem[6054] = 114;
razn_h_mem[6055] = 244;
razn_h_mem[6056] = 120;
razn_h_mem[6057] = 250;
razn_h_mem[6058] = 126;
razn_h_mem[6059] = 2;
razn_h_mem[6060] = 132;
razn_h_mem[6061] = 8;
razn_h_mem[6062] = 138;
razn_h_mem[6063] = 14;
razn_h_mem[6064] = 144;
razn_h_mem[6065] = 20;
razn_h_mem[6066] = 150;
razn_h_mem[6067] = 26;
razn_h_mem[6068] = 156;
razn_h_mem[6069] = 32;
razn_h_mem[6070] = 162;
razn_h_mem[6071] = 38;
razn_h_mem[6072] = 168;
razn_h_mem[6073] = 44;
razn_h_mem[6074] = 174;
razn_h_mem[6075] = 50;
razn_h_mem[6076] = 180;
razn_h_mem[6077] = 56;
razn_h_mem[6078] = 186;
razn_h_mem[6079] = 62;
razn_h_mem[6080] = 192;
razn_h_mem[6081] = 68;
razn_h_mem[6082] = 198;
razn_h_mem[6083] = 74;
razn_h_mem[6084] = 204;
razn_h_mem[6085] = 80;
razn_h_mem[6086] = 210;
razn_h_mem[6087] = 86;
razn_h_mem[6088] = 216;
razn_h_mem[6089] = 92;
razn_h_mem[6090] = 222;
razn_h_mem[6091] = 98;
razn_h_mem[6092] = 228;
razn_h_mem[6093] = 104;
razn_h_mem[6094] = 234;
razn_h_mem[6095] = 110;
razn_h_mem[6096] = 240;
razn_h_mem[6097] = 116;
razn_h_mem[6098] = 246;
razn_h_mem[6099] = 122;
razn_h_mem[6100] = 252;
razn_h_mem[6101] = 128;
razn_h_mem[6102] = 4;
razn_h_mem[6103] = 134;
razn_h_mem[6104] = 10;
razn_h_mem[6105] = 140;
razn_h_mem[6106] = 16;
razn_h_mem[6107] = 146;
razn_h_mem[6108] = 22;
razn_h_mem[6109] = 152;
razn_h_mem[6110] = 28;
razn_h_mem[6111] = 158;
razn_h_mem[6112] = 34;
razn_h_mem[6113] = 164;
razn_h_mem[6114] = 40;
razn_h_mem[6115] = 170;
razn_h_mem[6116] = 46;
razn_h_mem[6117] = 176;
razn_h_mem[6118] = 52;
razn_h_mem[6119] = 182;
razn_h_mem[6120] = 58;
razn_h_mem[6121] = 188;
razn_h_mem[6122] = 64;
razn_h_mem[6123] = 194;
razn_h_mem[6124] = 70;
razn_h_mem[6125] = 200;
razn_h_mem[6126] = 76;
razn_h_mem[6127] = 206;
razn_h_mem[6128] = 82;
razn_h_mem[6129] = 212;
razn_h_mem[6130] = 88;
razn_h_mem[6131] = 218;
razn_h_mem[6132] = 94;
razn_h_mem[6133] = 224;
razn_h_mem[6134] = 100;
razn_h_mem[6135] = 230;
razn_h_mem[6136] = 106;
razn_h_mem[6137] = 236;
razn_h_mem[6138] = 112;
razn_h_mem[6139] = 242;
razn_h_mem[6140] = 118;
razn_h_mem[6141] = 248;
razn_h_mem[6142] = 124;
razn_h_mem[6143] = 255;
razn_h_mem[6144] = 0;
razn_h_mem[6145] = 130;
razn_h_mem[6146] = 6;
razn_h_mem[6147] = 136;
razn_h_mem[6148] = 12;
razn_h_mem[6149] = 142;
razn_h_mem[6150] = 18;
razn_h_mem[6151] = 148;
razn_h_mem[6152] = 24;
razn_h_mem[6153] = 154;
razn_h_mem[6154] = 30;
razn_h_mem[6155] = 160;
razn_h_mem[6156] = 36;
razn_h_mem[6157] = 166;
razn_h_mem[6158] = 42;
razn_h_mem[6159] = 172;
razn_h_mem[6160] = 48;
razn_h_mem[6161] = 178;
razn_h_mem[6162] = 54;
razn_h_mem[6163] = 184;
razn_h_mem[6164] = 60;
razn_h_mem[6165] = 190;
razn_h_mem[6166] = 66;
razn_h_mem[6167] = 196;
razn_h_mem[6168] = 72;
razn_h_mem[6169] = 202;
razn_h_mem[6170] = 78;
razn_h_mem[6171] = 208;
razn_h_mem[6172] = 84;
razn_h_mem[6173] = 214;
razn_h_mem[6174] = 90;
razn_h_mem[6175] = 220;
razn_h_mem[6176] = 96;
razn_h_mem[6177] = 226;
razn_h_mem[6178] = 102;
razn_h_mem[6179] = 232;
razn_h_mem[6180] = 108;
razn_h_mem[6181] = 238;
razn_h_mem[6182] = 114;
razn_h_mem[6183] = 244;
razn_h_mem[6184] = 120;
razn_h_mem[6185] = 250;
razn_h_mem[6186] = 126;
razn_h_mem[6187] = 2;
razn_h_mem[6188] = 132;
razn_h_mem[6189] = 8;
razn_h_mem[6190] = 138;
razn_h_mem[6191] = 14;
razn_h_mem[6192] = 144;
razn_h_mem[6193] = 20;
razn_h_mem[6194] = 150;
razn_h_mem[6195] = 26;
razn_h_mem[6196] = 156;
razn_h_mem[6197] = 32;
razn_h_mem[6198] = 162;
razn_h_mem[6199] = 38;
razn_h_mem[6200] = 168;
razn_h_mem[6201] = 44;
razn_h_mem[6202] = 174;
razn_h_mem[6203] = 50;
razn_h_mem[6204] = 180;
razn_h_mem[6205] = 56;
razn_h_mem[6206] = 186;
razn_h_mem[6207] = 62;
razn_h_mem[6208] = 192;
razn_h_mem[6209] = 68;
razn_h_mem[6210] = 198;
razn_h_mem[6211] = 74;
razn_h_mem[6212] = 204;
razn_h_mem[6213] = 80;
razn_h_mem[6214] = 210;
razn_h_mem[6215] = 86;
razn_h_mem[6216] = 216;
razn_h_mem[6217] = 92;
razn_h_mem[6218] = 222;
razn_h_mem[6219] = 98;
razn_h_mem[6220] = 228;
razn_h_mem[6221] = 104;
razn_h_mem[6222] = 234;
razn_h_mem[6223] = 110;
razn_h_mem[6224] = 240;
razn_h_mem[6225] = 116;
razn_h_mem[6226] = 246;
razn_h_mem[6227] = 122;
razn_h_mem[6228] = 252;
razn_h_mem[6229] = 128;
razn_h_mem[6230] = 4;
razn_h_mem[6231] = 134;
razn_h_mem[6232] = 10;
razn_h_mem[6233] = 140;
razn_h_mem[6234] = 16;
razn_h_mem[6235] = 146;
razn_h_mem[6236] = 22;
razn_h_mem[6237] = 152;
razn_h_mem[6238] = 28;
razn_h_mem[6239] = 158;
razn_h_mem[6240] = 34;
razn_h_mem[6241] = 164;
razn_h_mem[6242] = 40;
razn_h_mem[6243] = 170;
razn_h_mem[6244] = 46;
razn_h_mem[6245] = 176;
razn_h_mem[6246] = 52;
razn_h_mem[6247] = 182;
razn_h_mem[6248] = 58;
razn_h_mem[6249] = 188;
razn_h_mem[6250] = 64;
razn_h_mem[6251] = 194;
razn_h_mem[6252] = 70;
razn_h_mem[6253] = 200;
razn_h_mem[6254] = 76;
razn_h_mem[6255] = 206;
razn_h_mem[6256] = 82;
razn_h_mem[6257] = 212;
razn_h_mem[6258] = 88;
razn_h_mem[6259] = 218;
razn_h_mem[6260] = 94;
razn_h_mem[6261] = 224;
razn_h_mem[6262] = 100;
razn_h_mem[6263] = 230;
razn_h_mem[6264] = 106;
razn_h_mem[6265] = 236;
razn_h_mem[6266] = 112;
razn_h_mem[6267] = 242;
razn_h_mem[6268] = 118;
razn_h_mem[6269] = 248;
razn_h_mem[6270] = 124;
razn_h_mem[6271] = 255;
razn_h_mem[6272] = 0;
razn_h_mem[6273] = 130;
razn_h_mem[6274] = 6;
razn_h_mem[6275] = 136;
razn_h_mem[6276] = 12;
razn_h_mem[6277] = 142;
razn_h_mem[6278] = 18;
razn_h_mem[6279] = 148;
razn_h_mem[6280] = 24;
razn_h_mem[6281] = 154;
razn_h_mem[6282] = 30;
razn_h_mem[6283] = 160;
razn_h_mem[6284] = 36;
razn_h_mem[6285] = 166;
razn_h_mem[6286] = 42;
razn_h_mem[6287] = 172;
razn_h_mem[6288] = 48;
razn_h_mem[6289] = 178;
razn_h_mem[6290] = 54;
razn_h_mem[6291] = 184;
razn_h_mem[6292] = 60;
razn_h_mem[6293] = 190;
razn_h_mem[6294] = 66;
razn_h_mem[6295] = 196;
razn_h_mem[6296] = 72;
razn_h_mem[6297] = 202;
razn_h_mem[6298] = 78;
razn_h_mem[6299] = 208;
razn_h_mem[6300] = 84;
razn_h_mem[6301] = 214;
razn_h_mem[6302] = 90;
razn_h_mem[6303] = 220;
razn_h_mem[6304] = 96;
razn_h_mem[6305] = 226;
razn_h_mem[6306] = 102;
razn_h_mem[6307] = 232;
razn_h_mem[6308] = 108;
razn_h_mem[6309] = 238;
razn_h_mem[6310] = 114;
razn_h_mem[6311] = 244;
razn_h_mem[6312] = 120;
razn_h_mem[6313] = 250;
razn_h_mem[6314] = 126;
razn_h_mem[6315] = 2;
razn_h_mem[6316] = 132;
razn_h_mem[6317] = 8;
razn_h_mem[6318] = 138;
razn_h_mem[6319] = 14;
razn_h_mem[6320] = 144;
razn_h_mem[6321] = 20;
razn_h_mem[6322] = 150;
razn_h_mem[6323] = 26;
razn_h_mem[6324] = 156;
razn_h_mem[6325] = 32;
razn_h_mem[6326] = 162;
razn_h_mem[6327] = 38;
razn_h_mem[6328] = 168;
razn_h_mem[6329] = 44;
razn_h_mem[6330] = 174;
razn_h_mem[6331] = 50;
razn_h_mem[6332] = 180;
razn_h_mem[6333] = 56;
razn_h_mem[6334] = 186;
razn_h_mem[6335] = 62;
razn_h_mem[6336] = 192;
razn_h_mem[6337] = 68;
razn_h_mem[6338] = 198;
razn_h_mem[6339] = 74;
razn_h_mem[6340] = 204;
razn_h_mem[6341] = 80;
razn_h_mem[6342] = 210;
razn_h_mem[6343] = 86;
razn_h_mem[6344] = 216;
razn_h_mem[6345] = 92;
razn_h_mem[6346] = 222;
razn_h_mem[6347] = 98;
razn_h_mem[6348] = 228;
razn_h_mem[6349] = 104;
razn_h_mem[6350] = 234;
razn_h_mem[6351] = 110;
razn_h_mem[6352] = 240;
razn_h_mem[6353] = 116;
razn_h_mem[6354] = 246;
razn_h_mem[6355] = 122;
razn_h_mem[6356] = 252;
razn_h_mem[6357] = 128;
razn_h_mem[6358] = 4;
razn_h_mem[6359] = 134;
razn_h_mem[6360] = 10;
razn_h_mem[6361] = 140;
razn_h_mem[6362] = 16;
razn_h_mem[6363] = 146;
razn_h_mem[6364] = 22;
razn_h_mem[6365] = 152;
razn_h_mem[6366] = 28;
razn_h_mem[6367] = 158;
razn_h_mem[6368] = 34;
razn_h_mem[6369] = 164;
razn_h_mem[6370] = 40;
razn_h_mem[6371] = 170;
razn_h_mem[6372] = 46;
razn_h_mem[6373] = 176;
razn_h_mem[6374] = 52;
razn_h_mem[6375] = 182;
razn_h_mem[6376] = 58;
razn_h_mem[6377] = 188;
razn_h_mem[6378] = 64;
razn_h_mem[6379] = 194;
razn_h_mem[6380] = 70;
razn_h_mem[6381] = 200;
razn_h_mem[6382] = 76;
razn_h_mem[6383] = 206;
razn_h_mem[6384] = 82;
razn_h_mem[6385] = 212;
razn_h_mem[6386] = 88;
razn_h_mem[6387] = 218;
razn_h_mem[6388] = 94;
razn_h_mem[6389] = 224;
razn_h_mem[6390] = 100;
razn_h_mem[6391] = 230;
razn_h_mem[6392] = 106;
razn_h_mem[6393] = 236;
razn_h_mem[6394] = 112;
razn_h_mem[6395] = 242;
razn_h_mem[6396] = 118;
razn_h_mem[6397] = 248;
razn_h_mem[6398] = 124;
razn_h_mem[6399] = 255;
razn_h_mem[6400] = 0;
razn_h_mem[6401] = 130;
razn_h_mem[6402] = 6;
razn_h_mem[6403] = 136;
razn_h_mem[6404] = 12;
razn_h_mem[6405] = 142;
razn_h_mem[6406] = 18;
razn_h_mem[6407] = 148;
razn_h_mem[6408] = 24;
razn_h_mem[6409] = 154;
razn_h_mem[6410] = 30;
razn_h_mem[6411] = 160;
razn_h_mem[6412] = 36;
razn_h_mem[6413] = 166;
razn_h_mem[6414] = 42;
razn_h_mem[6415] = 172;
razn_h_mem[6416] = 48;
razn_h_mem[6417] = 178;
razn_h_mem[6418] = 54;
razn_h_mem[6419] = 184;
razn_h_mem[6420] = 60;
razn_h_mem[6421] = 190;
razn_h_mem[6422] = 66;
razn_h_mem[6423] = 196;
razn_h_mem[6424] = 72;
razn_h_mem[6425] = 202;
razn_h_mem[6426] = 78;
razn_h_mem[6427] = 208;
razn_h_mem[6428] = 84;
razn_h_mem[6429] = 214;
razn_h_mem[6430] = 90;
razn_h_mem[6431] = 220;
razn_h_mem[6432] = 96;
razn_h_mem[6433] = 226;
razn_h_mem[6434] = 102;
razn_h_mem[6435] = 232;
razn_h_mem[6436] = 108;
razn_h_mem[6437] = 238;
razn_h_mem[6438] = 114;
razn_h_mem[6439] = 244;
razn_h_mem[6440] = 120;
razn_h_mem[6441] = 250;
razn_h_mem[6442] = 126;
razn_h_mem[6443] = 2;
razn_h_mem[6444] = 132;
razn_h_mem[6445] = 8;
razn_h_mem[6446] = 138;
razn_h_mem[6447] = 14;
razn_h_mem[6448] = 144;
razn_h_mem[6449] = 20;
razn_h_mem[6450] = 150;
razn_h_mem[6451] = 26;
razn_h_mem[6452] = 156;
razn_h_mem[6453] = 32;
razn_h_mem[6454] = 162;
razn_h_mem[6455] = 38;
razn_h_mem[6456] = 168;
razn_h_mem[6457] = 44;
razn_h_mem[6458] = 174;
razn_h_mem[6459] = 50;
razn_h_mem[6460] = 180;
razn_h_mem[6461] = 56;
razn_h_mem[6462] = 186;
razn_h_mem[6463] = 62;
razn_h_mem[6464] = 192;
razn_h_mem[6465] = 68;
razn_h_mem[6466] = 198;
razn_h_mem[6467] = 74;
razn_h_mem[6468] = 204;
razn_h_mem[6469] = 80;
razn_h_mem[6470] = 210;
razn_h_mem[6471] = 86;
razn_h_mem[6472] = 216;
razn_h_mem[6473] = 92;
razn_h_mem[6474] = 222;
razn_h_mem[6475] = 98;
razn_h_mem[6476] = 228;
razn_h_mem[6477] = 104;
razn_h_mem[6478] = 234;
razn_h_mem[6479] = 110;
razn_h_mem[6480] = 240;
razn_h_mem[6481] = 116;
razn_h_mem[6482] = 246;
razn_h_mem[6483] = 122;
razn_h_mem[6484] = 252;
razn_h_mem[6485] = 128;
razn_h_mem[6486] = 4;
razn_h_mem[6487] = 134;
razn_h_mem[6488] = 10;
razn_h_mem[6489] = 140;
razn_h_mem[6490] = 16;
razn_h_mem[6491] = 146;
razn_h_mem[6492] = 22;
razn_h_mem[6493] = 152;
razn_h_mem[6494] = 28;
razn_h_mem[6495] = 158;
razn_h_mem[6496] = 34;
razn_h_mem[6497] = 164;
razn_h_mem[6498] = 40;
razn_h_mem[6499] = 170;
razn_h_mem[6500] = 46;
razn_h_mem[6501] = 176;
razn_h_mem[6502] = 52;
razn_h_mem[6503] = 182;
razn_h_mem[6504] = 58;
razn_h_mem[6505] = 188;
razn_h_mem[6506] = 64;
razn_h_mem[6507] = 194;
razn_h_mem[6508] = 70;
razn_h_mem[6509] = 200;
razn_h_mem[6510] = 76;
razn_h_mem[6511] = 206;
razn_h_mem[6512] = 82;
razn_h_mem[6513] = 212;
razn_h_mem[6514] = 88;
razn_h_mem[6515] = 218;
razn_h_mem[6516] = 94;
razn_h_mem[6517] = 224;
razn_h_mem[6518] = 100;
razn_h_mem[6519] = 230;
razn_h_mem[6520] = 106;
razn_h_mem[6521] = 236;
razn_h_mem[6522] = 112;
razn_h_mem[6523] = 242;
razn_h_mem[6524] = 118;
razn_h_mem[6525] = 248;
razn_h_mem[6526] = 124;
razn_h_mem[6527] = 255;
razn_h_mem[6528] = 0;
razn_h_mem[6529] = 130;
razn_h_mem[6530] = 6;
razn_h_mem[6531] = 136;
razn_h_mem[6532] = 12;
razn_h_mem[6533] = 142;
razn_h_mem[6534] = 18;
razn_h_mem[6535] = 148;
razn_h_mem[6536] = 24;
razn_h_mem[6537] = 154;
razn_h_mem[6538] = 30;
razn_h_mem[6539] = 160;
razn_h_mem[6540] = 36;
razn_h_mem[6541] = 166;
razn_h_mem[6542] = 42;
razn_h_mem[6543] = 172;
razn_h_mem[6544] = 48;
razn_h_mem[6545] = 178;
razn_h_mem[6546] = 54;
razn_h_mem[6547] = 184;
razn_h_mem[6548] = 60;
razn_h_mem[6549] = 190;
razn_h_mem[6550] = 66;
razn_h_mem[6551] = 196;
razn_h_mem[6552] = 72;
razn_h_mem[6553] = 202;
razn_h_mem[6554] = 78;
razn_h_mem[6555] = 208;
razn_h_mem[6556] = 84;
razn_h_mem[6557] = 214;
razn_h_mem[6558] = 90;
razn_h_mem[6559] = 220;
razn_h_mem[6560] = 96;
razn_h_mem[6561] = 226;
razn_h_mem[6562] = 102;
razn_h_mem[6563] = 232;
razn_h_mem[6564] = 108;
razn_h_mem[6565] = 238;
razn_h_mem[6566] = 114;
razn_h_mem[6567] = 244;
razn_h_mem[6568] = 120;
razn_h_mem[6569] = 250;
razn_h_mem[6570] = 126;
razn_h_mem[6571] = 2;
razn_h_mem[6572] = 132;
razn_h_mem[6573] = 8;
razn_h_mem[6574] = 138;
razn_h_mem[6575] = 14;
razn_h_mem[6576] = 144;
razn_h_mem[6577] = 20;
razn_h_mem[6578] = 150;
razn_h_mem[6579] = 26;
razn_h_mem[6580] = 156;
razn_h_mem[6581] = 32;
razn_h_mem[6582] = 162;
razn_h_mem[6583] = 38;
razn_h_mem[6584] = 168;
razn_h_mem[6585] = 44;
razn_h_mem[6586] = 174;
razn_h_mem[6587] = 50;
razn_h_mem[6588] = 180;
razn_h_mem[6589] = 56;
razn_h_mem[6590] = 186;
razn_h_mem[6591] = 62;
razn_h_mem[6592] = 192;
razn_h_mem[6593] = 68;
razn_h_mem[6594] = 198;
razn_h_mem[6595] = 74;
razn_h_mem[6596] = 204;
razn_h_mem[6597] = 80;
razn_h_mem[6598] = 210;
razn_h_mem[6599] = 86;
razn_h_mem[6600] = 216;
razn_h_mem[6601] = 92;
razn_h_mem[6602] = 222;
razn_h_mem[6603] = 98;
razn_h_mem[6604] = 228;
razn_h_mem[6605] = 104;
razn_h_mem[6606] = 234;
razn_h_mem[6607] = 110;
razn_h_mem[6608] = 240;
razn_h_mem[6609] = 116;
razn_h_mem[6610] = 246;
razn_h_mem[6611] = 122;
razn_h_mem[6612] = 252;
razn_h_mem[6613] = 128;
razn_h_mem[6614] = 4;
razn_h_mem[6615] = 134;
razn_h_mem[6616] = 10;
razn_h_mem[6617] = 140;
razn_h_mem[6618] = 16;
razn_h_mem[6619] = 146;
razn_h_mem[6620] = 22;
razn_h_mem[6621] = 152;
razn_h_mem[6622] = 28;
razn_h_mem[6623] = 158;
razn_h_mem[6624] = 34;
razn_h_mem[6625] = 164;
razn_h_mem[6626] = 40;
razn_h_mem[6627] = 170;
razn_h_mem[6628] = 46;
razn_h_mem[6629] = 176;
razn_h_mem[6630] = 52;
razn_h_mem[6631] = 182;
razn_h_mem[6632] = 58;
razn_h_mem[6633] = 188;
razn_h_mem[6634] = 64;
razn_h_mem[6635] = 194;
razn_h_mem[6636] = 70;
razn_h_mem[6637] = 200;
razn_h_mem[6638] = 76;
razn_h_mem[6639] = 206;
razn_h_mem[6640] = 82;
razn_h_mem[6641] = 212;
razn_h_mem[6642] = 88;
razn_h_mem[6643] = 218;
razn_h_mem[6644] = 94;
razn_h_mem[6645] = 224;
razn_h_mem[6646] = 100;
razn_h_mem[6647] = 230;
razn_h_mem[6648] = 106;
razn_h_mem[6649] = 236;
razn_h_mem[6650] = 112;
razn_h_mem[6651] = 242;
razn_h_mem[6652] = 118;
razn_h_mem[6653] = 248;
razn_h_mem[6654] = 124;
razn_h_mem[6655] = 255;
razn_h_mem[6656] = 0;
razn_h_mem[6657] = 130;
razn_h_mem[6658] = 6;
razn_h_mem[6659] = 136;
razn_h_mem[6660] = 12;
razn_h_mem[6661] = 142;
razn_h_mem[6662] = 18;
razn_h_mem[6663] = 148;
razn_h_mem[6664] = 24;
razn_h_mem[6665] = 154;
razn_h_mem[6666] = 30;
razn_h_mem[6667] = 160;
razn_h_mem[6668] = 36;
razn_h_mem[6669] = 166;
razn_h_mem[6670] = 42;
razn_h_mem[6671] = 172;
razn_h_mem[6672] = 48;
razn_h_mem[6673] = 178;
razn_h_mem[6674] = 54;
razn_h_mem[6675] = 184;
razn_h_mem[6676] = 60;
razn_h_mem[6677] = 190;
razn_h_mem[6678] = 66;
razn_h_mem[6679] = 196;
razn_h_mem[6680] = 72;
razn_h_mem[6681] = 202;
razn_h_mem[6682] = 78;
razn_h_mem[6683] = 208;
razn_h_mem[6684] = 84;
razn_h_mem[6685] = 214;
razn_h_mem[6686] = 90;
razn_h_mem[6687] = 220;
razn_h_mem[6688] = 96;
razn_h_mem[6689] = 226;
razn_h_mem[6690] = 102;
razn_h_mem[6691] = 232;
razn_h_mem[6692] = 108;
razn_h_mem[6693] = 238;
razn_h_mem[6694] = 114;
razn_h_mem[6695] = 244;
razn_h_mem[6696] = 120;
razn_h_mem[6697] = 250;
razn_h_mem[6698] = 126;
razn_h_mem[6699] = 2;
razn_h_mem[6700] = 132;
razn_h_mem[6701] = 8;
razn_h_mem[6702] = 138;
razn_h_mem[6703] = 14;
razn_h_mem[6704] = 144;
razn_h_mem[6705] = 20;
razn_h_mem[6706] = 150;
razn_h_mem[6707] = 26;
razn_h_mem[6708] = 156;
razn_h_mem[6709] = 32;
razn_h_mem[6710] = 162;
razn_h_mem[6711] = 38;
razn_h_mem[6712] = 168;
razn_h_mem[6713] = 44;
razn_h_mem[6714] = 174;
razn_h_mem[6715] = 50;
razn_h_mem[6716] = 180;
razn_h_mem[6717] = 56;
razn_h_mem[6718] = 186;
razn_h_mem[6719] = 62;
razn_h_mem[6720] = 192;
razn_h_mem[6721] = 68;
razn_h_mem[6722] = 198;
razn_h_mem[6723] = 74;
razn_h_mem[6724] = 204;
razn_h_mem[6725] = 80;
razn_h_mem[6726] = 210;
razn_h_mem[6727] = 86;
razn_h_mem[6728] = 216;
razn_h_mem[6729] = 92;
razn_h_mem[6730] = 222;
razn_h_mem[6731] = 98;
razn_h_mem[6732] = 228;
razn_h_mem[6733] = 104;
razn_h_mem[6734] = 234;
razn_h_mem[6735] = 110;
razn_h_mem[6736] = 240;
razn_h_mem[6737] = 116;
razn_h_mem[6738] = 246;
razn_h_mem[6739] = 122;
razn_h_mem[6740] = 252;
razn_h_mem[6741] = 128;
razn_h_mem[6742] = 4;
razn_h_mem[6743] = 134;
razn_h_mem[6744] = 10;
razn_h_mem[6745] = 140;
razn_h_mem[6746] = 16;
razn_h_mem[6747] = 146;
razn_h_mem[6748] = 22;
razn_h_mem[6749] = 152;
razn_h_mem[6750] = 28;
razn_h_mem[6751] = 158;
razn_h_mem[6752] = 34;
razn_h_mem[6753] = 164;
razn_h_mem[6754] = 40;
razn_h_mem[6755] = 170;
razn_h_mem[6756] = 46;
razn_h_mem[6757] = 176;
razn_h_mem[6758] = 52;
razn_h_mem[6759] = 182;
razn_h_mem[6760] = 58;
razn_h_mem[6761] = 188;
razn_h_mem[6762] = 64;
razn_h_mem[6763] = 194;
razn_h_mem[6764] = 70;
razn_h_mem[6765] = 200;
razn_h_mem[6766] = 76;
razn_h_mem[6767] = 206;
razn_h_mem[6768] = 82;
razn_h_mem[6769] = 212;
razn_h_mem[6770] = 88;
razn_h_mem[6771] = 218;
razn_h_mem[6772] = 94;
razn_h_mem[6773] = 224;
razn_h_mem[6774] = 100;
razn_h_mem[6775] = 230;
razn_h_mem[6776] = 106;
razn_h_mem[6777] = 236;
razn_h_mem[6778] = 112;
razn_h_mem[6779] = 242;
razn_h_mem[6780] = 118;
razn_h_mem[6781] = 248;
razn_h_mem[6782] = 124;
razn_h_mem[6783] = 255;
razn_h_mem[6784] = 0;
razn_h_mem[6785] = 130;
razn_h_mem[6786] = 6;
razn_h_mem[6787] = 136;
razn_h_mem[6788] = 12;
razn_h_mem[6789] = 142;
razn_h_mem[6790] = 18;
razn_h_mem[6791] = 148;
razn_h_mem[6792] = 24;
razn_h_mem[6793] = 154;
razn_h_mem[6794] = 30;
razn_h_mem[6795] = 160;
razn_h_mem[6796] = 36;
razn_h_mem[6797] = 166;
razn_h_mem[6798] = 42;
razn_h_mem[6799] = 172;
razn_h_mem[6800] = 48;
razn_h_mem[6801] = 178;
razn_h_mem[6802] = 54;
razn_h_mem[6803] = 184;
razn_h_mem[6804] = 60;
razn_h_mem[6805] = 190;
razn_h_mem[6806] = 66;
razn_h_mem[6807] = 196;
razn_h_mem[6808] = 72;
razn_h_mem[6809] = 202;
razn_h_mem[6810] = 78;
razn_h_mem[6811] = 208;
razn_h_mem[6812] = 84;
razn_h_mem[6813] = 214;
razn_h_mem[6814] = 90;
razn_h_mem[6815] = 220;
razn_h_mem[6816] = 96;
razn_h_mem[6817] = 226;
razn_h_mem[6818] = 102;
razn_h_mem[6819] = 232;
razn_h_mem[6820] = 108;
razn_h_mem[6821] = 238;
razn_h_mem[6822] = 114;
razn_h_mem[6823] = 244;
razn_h_mem[6824] = 120;
razn_h_mem[6825] = 250;
razn_h_mem[6826] = 126;
razn_h_mem[6827] = 2;
razn_h_mem[6828] = 132;
razn_h_mem[6829] = 8;
razn_h_mem[6830] = 138;
razn_h_mem[6831] = 14;
razn_h_mem[6832] = 144;
razn_h_mem[6833] = 20;
razn_h_mem[6834] = 150;
razn_h_mem[6835] = 26;
razn_h_mem[6836] = 156;
razn_h_mem[6837] = 32;
razn_h_mem[6838] = 162;
razn_h_mem[6839] = 38;
razn_h_mem[6840] = 168;
razn_h_mem[6841] = 44;
razn_h_mem[6842] = 174;
razn_h_mem[6843] = 50;
razn_h_mem[6844] = 180;
razn_h_mem[6845] = 56;
razn_h_mem[6846] = 186;
razn_h_mem[6847] = 62;
razn_h_mem[6848] = 192;
razn_h_mem[6849] = 68;
razn_h_mem[6850] = 198;
razn_h_mem[6851] = 74;
razn_h_mem[6852] = 204;
razn_h_mem[6853] = 80;
razn_h_mem[6854] = 210;
razn_h_mem[6855] = 86;
razn_h_mem[6856] = 216;
razn_h_mem[6857] = 92;
razn_h_mem[6858] = 222;
razn_h_mem[6859] = 98;
razn_h_mem[6860] = 228;
razn_h_mem[6861] = 104;
razn_h_mem[6862] = 234;
razn_h_mem[6863] = 110;
razn_h_mem[6864] = 240;
razn_h_mem[6865] = 116;
razn_h_mem[6866] = 246;
razn_h_mem[6867] = 122;
razn_h_mem[6868] = 252;
razn_h_mem[6869] = 128;
razn_h_mem[6870] = 4;
razn_h_mem[6871] = 134;
razn_h_mem[6872] = 10;
razn_h_mem[6873] = 140;
razn_h_mem[6874] = 16;
razn_h_mem[6875] = 146;
razn_h_mem[6876] = 22;
razn_h_mem[6877] = 152;
razn_h_mem[6878] = 28;
razn_h_mem[6879] = 158;
razn_h_mem[6880] = 34;
razn_h_mem[6881] = 164;
razn_h_mem[6882] = 40;
razn_h_mem[6883] = 170;
razn_h_mem[6884] = 46;
razn_h_mem[6885] = 176;
razn_h_mem[6886] = 52;
razn_h_mem[6887] = 182;
razn_h_mem[6888] = 58;
razn_h_mem[6889] = 188;
razn_h_mem[6890] = 64;
razn_h_mem[6891] = 194;
razn_h_mem[6892] = 70;
razn_h_mem[6893] = 200;
razn_h_mem[6894] = 76;
razn_h_mem[6895] = 206;
razn_h_mem[6896] = 82;
razn_h_mem[6897] = 212;
razn_h_mem[6898] = 88;
razn_h_mem[6899] = 218;
razn_h_mem[6900] = 94;
razn_h_mem[6901] = 224;
razn_h_mem[6902] = 100;
razn_h_mem[6903] = 230;
razn_h_mem[6904] = 106;
razn_h_mem[6905] = 236;
razn_h_mem[6906] = 112;
razn_h_mem[6907] = 242;
razn_h_mem[6908] = 118;
razn_h_mem[6909] = 248;
razn_h_mem[6910] = 124;
razn_h_mem[6911] = 255;
razn_h_mem[6912] = 0;
razn_h_mem[6913] = 130;
razn_h_mem[6914] = 6;
razn_h_mem[6915] = 136;
razn_h_mem[6916] = 12;
razn_h_mem[6917] = 142;
razn_h_mem[6918] = 18;
razn_h_mem[6919] = 148;
razn_h_mem[6920] = 24;
razn_h_mem[6921] = 154;
razn_h_mem[6922] = 30;
razn_h_mem[6923] = 160;
razn_h_mem[6924] = 36;
razn_h_mem[6925] = 166;
razn_h_mem[6926] = 42;
razn_h_mem[6927] = 172;
razn_h_mem[6928] = 48;
razn_h_mem[6929] = 178;
razn_h_mem[6930] = 54;
razn_h_mem[6931] = 184;
razn_h_mem[6932] = 60;
razn_h_mem[6933] = 190;
razn_h_mem[6934] = 66;
razn_h_mem[6935] = 196;
razn_h_mem[6936] = 72;
razn_h_mem[6937] = 202;
razn_h_mem[6938] = 78;
razn_h_mem[6939] = 208;
razn_h_mem[6940] = 84;
razn_h_mem[6941] = 214;
razn_h_mem[6942] = 90;
razn_h_mem[6943] = 220;
razn_h_mem[6944] = 96;
razn_h_mem[6945] = 226;
razn_h_mem[6946] = 102;
razn_h_mem[6947] = 232;
razn_h_mem[6948] = 108;
razn_h_mem[6949] = 238;
razn_h_mem[6950] = 114;
razn_h_mem[6951] = 244;
razn_h_mem[6952] = 120;
razn_h_mem[6953] = 250;
razn_h_mem[6954] = 126;
razn_h_mem[6955] = 2;
razn_h_mem[6956] = 132;
razn_h_mem[6957] = 8;
razn_h_mem[6958] = 138;
razn_h_mem[6959] = 14;
razn_h_mem[6960] = 144;
razn_h_mem[6961] = 20;
razn_h_mem[6962] = 150;
razn_h_mem[6963] = 26;
razn_h_mem[6964] = 156;
razn_h_mem[6965] = 32;
razn_h_mem[6966] = 162;
razn_h_mem[6967] = 38;
razn_h_mem[6968] = 168;
razn_h_mem[6969] = 44;
razn_h_mem[6970] = 174;
razn_h_mem[6971] = 50;
razn_h_mem[6972] = 180;
razn_h_mem[6973] = 56;
razn_h_mem[6974] = 186;
razn_h_mem[6975] = 62;
razn_h_mem[6976] = 192;
razn_h_mem[6977] = 68;
razn_h_mem[6978] = 198;
razn_h_mem[6979] = 74;
razn_h_mem[6980] = 204;
razn_h_mem[6981] = 80;
razn_h_mem[6982] = 210;
razn_h_mem[6983] = 86;
razn_h_mem[6984] = 216;
razn_h_mem[6985] = 92;
razn_h_mem[6986] = 222;
razn_h_mem[6987] = 98;
razn_h_mem[6988] = 228;
razn_h_mem[6989] = 104;
razn_h_mem[6990] = 234;
razn_h_mem[6991] = 110;
razn_h_mem[6992] = 240;
razn_h_mem[6993] = 116;
razn_h_mem[6994] = 246;
razn_h_mem[6995] = 122;
razn_h_mem[6996] = 252;
razn_h_mem[6997] = 128;
razn_h_mem[6998] = 4;
razn_h_mem[6999] = 134;
razn_h_mem[7000] = 10;
razn_h_mem[7001] = 140;
razn_h_mem[7002] = 16;
razn_h_mem[7003] = 146;
razn_h_mem[7004] = 22;
razn_h_mem[7005] = 152;
razn_h_mem[7006] = 28;
razn_h_mem[7007] = 158;
razn_h_mem[7008] = 34;
razn_h_mem[7009] = 164;
razn_h_mem[7010] = 40;
razn_h_mem[7011] = 170;
razn_h_mem[7012] = 46;
razn_h_mem[7013] = 176;
razn_h_mem[7014] = 52;
razn_h_mem[7015] = 182;
razn_h_mem[7016] = 58;
razn_h_mem[7017] = 188;
razn_h_mem[7018] = 64;
razn_h_mem[7019] = 194;
razn_h_mem[7020] = 70;
razn_h_mem[7021] = 200;
razn_h_mem[7022] = 76;
razn_h_mem[7023] = 206;
razn_h_mem[7024] = 82;
razn_h_mem[7025] = 212;
razn_h_mem[7026] = 88;
razn_h_mem[7027] = 218;
razn_h_mem[7028] = 94;
razn_h_mem[7029] = 224;
razn_h_mem[7030] = 100;
razn_h_mem[7031] = 230;
razn_h_mem[7032] = 106;
razn_h_mem[7033] = 236;
razn_h_mem[7034] = 112;
razn_h_mem[7035] = 242;
razn_h_mem[7036] = 118;
razn_h_mem[7037] = 248;
razn_h_mem[7038] = 124;
razn_h_mem[7039] = 255;
razn_h_mem[7040] = 0;
razn_h_mem[7041] = 130;
razn_h_mem[7042] = 6;
razn_h_mem[7043] = 136;
razn_h_mem[7044] = 12;
razn_h_mem[7045] = 142;
razn_h_mem[7046] = 18;
razn_h_mem[7047] = 148;
razn_h_mem[7048] = 24;
razn_h_mem[7049] = 154;
razn_h_mem[7050] = 30;
razn_h_mem[7051] = 160;
razn_h_mem[7052] = 36;
razn_h_mem[7053] = 166;
razn_h_mem[7054] = 42;
razn_h_mem[7055] = 172;
razn_h_mem[7056] = 48;
razn_h_mem[7057] = 178;
razn_h_mem[7058] = 54;
razn_h_mem[7059] = 184;
razn_h_mem[7060] = 60;
razn_h_mem[7061] = 190;
razn_h_mem[7062] = 66;
razn_h_mem[7063] = 196;
razn_h_mem[7064] = 72;
razn_h_mem[7065] = 202;
razn_h_mem[7066] = 78;
razn_h_mem[7067] = 208;
razn_h_mem[7068] = 84;
razn_h_mem[7069] = 214;
razn_h_mem[7070] = 90;
razn_h_mem[7071] = 220;
razn_h_mem[7072] = 96;
razn_h_mem[7073] = 226;
razn_h_mem[7074] = 102;
razn_h_mem[7075] = 232;
razn_h_mem[7076] = 108;
razn_h_mem[7077] = 238;
razn_h_mem[7078] = 114;
razn_h_mem[7079] = 244;
razn_h_mem[7080] = 120;
razn_h_mem[7081] = 250;
razn_h_mem[7082] = 126;
razn_h_mem[7083] = 2;
razn_h_mem[7084] = 132;
razn_h_mem[7085] = 8;
razn_h_mem[7086] = 138;
razn_h_mem[7087] = 14;
razn_h_mem[7088] = 144;
razn_h_mem[7089] = 20;
razn_h_mem[7090] = 150;
razn_h_mem[7091] = 26;
razn_h_mem[7092] = 156;
razn_h_mem[7093] = 32;
razn_h_mem[7094] = 162;
razn_h_mem[7095] = 38;
razn_h_mem[7096] = 168;
razn_h_mem[7097] = 44;
razn_h_mem[7098] = 174;
razn_h_mem[7099] = 50;
razn_h_mem[7100] = 180;
razn_h_mem[7101] = 56;
razn_h_mem[7102] = 186;
razn_h_mem[7103] = 62;
razn_h_mem[7104] = 192;
razn_h_mem[7105] = 68;
razn_h_mem[7106] = 198;
razn_h_mem[7107] = 74;
razn_h_mem[7108] = 204;
razn_h_mem[7109] = 80;
razn_h_mem[7110] = 210;
razn_h_mem[7111] = 86;
razn_h_mem[7112] = 216;
razn_h_mem[7113] = 92;
razn_h_mem[7114] = 222;
razn_h_mem[7115] = 98;
razn_h_mem[7116] = 228;
razn_h_mem[7117] = 104;
razn_h_mem[7118] = 234;
razn_h_mem[7119] = 110;
razn_h_mem[7120] = 240;
razn_h_mem[7121] = 116;
razn_h_mem[7122] = 246;
razn_h_mem[7123] = 122;
razn_h_mem[7124] = 252;
razn_h_mem[7125] = 128;
razn_h_mem[7126] = 4;
razn_h_mem[7127] = 134;
razn_h_mem[7128] = 10;
razn_h_mem[7129] = 140;
razn_h_mem[7130] = 16;
razn_h_mem[7131] = 146;
razn_h_mem[7132] = 22;
razn_h_mem[7133] = 152;
razn_h_mem[7134] = 28;
razn_h_mem[7135] = 158;
razn_h_mem[7136] = 34;
razn_h_mem[7137] = 164;
razn_h_mem[7138] = 40;
razn_h_mem[7139] = 170;
razn_h_mem[7140] = 46;
razn_h_mem[7141] = 176;
razn_h_mem[7142] = 52;
razn_h_mem[7143] = 182;
razn_h_mem[7144] = 58;
razn_h_mem[7145] = 188;
razn_h_mem[7146] = 64;
razn_h_mem[7147] = 194;
razn_h_mem[7148] = 70;
razn_h_mem[7149] = 200;
razn_h_mem[7150] = 76;
razn_h_mem[7151] = 206;
razn_h_mem[7152] = 82;
razn_h_mem[7153] = 212;
razn_h_mem[7154] = 88;
razn_h_mem[7155] = 218;
razn_h_mem[7156] = 94;
razn_h_mem[7157] = 224;
razn_h_mem[7158] = 100;
razn_h_mem[7159] = 230;
razn_h_mem[7160] = 106;
razn_h_mem[7161] = 236;
razn_h_mem[7162] = 112;
razn_h_mem[7163] = 242;
razn_h_mem[7164] = 118;
razn_h_mem[7165] = 248;
razn_h_mem[7166] = 124;
razn_h_mem[7167] = 255;
razn_h_mem[7168] = 0;
razn_h_mem[7169] = 130;
razn_h_mem[7170] = 6;
razn_h_mem[7171] = 136;
razn_h_mem[7172] = 12;
razn_h_mem[7173] = 142;
razn_h_mem[7174] = 18;
razn_h_mem[7175] = 148;
razn_h_mem[7176] = 24;
razn_h_mem[7177] = 154;
razn_h_mem[7178] = 30;
razn_h_mem[7179] = 160;
razn_h_mem[7180] = 36;
razn_h_mem[7181] = 166;
razn_h_mem[7182] = 42;
razn_h_mem[7183] = 172;
razn_h_mem[7184] = 48;
razn_h_mem[7185] = 178;
razn_h_mem[7186] = 54;
razn_h_mem[7187] = 184;
razn_h_mem[7188] = 60;
razn_h_mem[7189] = 190;
razn_h_mem[7190] = 66;
razn_h_mem[7191] = 196;
razn_h_mem[7192] = 72;
razn_h_mem[7193] = 202;
razn_h_mem[7194] = 78;
razn_h_mem[7195] = 208;
razn_h_mem[7196] = 84;
razn_h_mem[7197] = 214;
razn_h_mem[7198] = 90;
razn_h_mem[7199] = 220;
razn_h_mem[7200] = 96;
razn_h_mem[7201] = 226;
razn_h_mem[7202] = 102;
razn_h_mem[7203] = 232;
razn_h_mem[7204] = 108;
razn_h_mem[7205] = 238;
razn_h_mem[7206] = 114;
razn_h_mem[7207] = 244;
razn_h_mem[7208] = 120;
razn_h_mem[7209] = 250;
razn_h_mem[7210] = 126;
razn_h_mem[7211] = 2;
razn_h_mem[7212] = 132;
razn_h_mem[7213] = 8;
razn_h_mem[7214] = 138;
razn_h_mem[7215] = 14;
razn_h_mem[7216] = 144;
razn_h_mem[7217] = 20;
razn_h_mem[7218] = 150;
razn_h_mem[7219] = 26;
razn_h_mem[7220] = 156;
razn_h_mem[7221] = 32;
razn_h_mem[7222] = 162;
razn_h_mem[7223] = 38;
razn_h_mem[7224] = 168;
razn_h_mem[7225] = 44;
razn_h_mem[7226] = 174;
razn_h_mem[7227] = 50;
razn_h_mem[7228] = 180;
razn_h_mem[7229] = 56;
razn_h_mem[7230] = 186;
razn_h_mem[7231] = 62;
razn_h_mem[7232] = 192;
razn_h_mem[7233] = 68;
razn_h_mem[7234] = 198;
razn_h_mem[7235] = 74;
razn_h_mem[7236] = 204;
razn_h_mem[7237] = 80;
razn_h_mem[7238] = 210;
razn_h_mem[7239] = 86;
razn_h_mem[7240] = 216;
razn_h_mem[7241] = 92;
razn_h_mem[7242] = 222;
razn_h_mem[7243] = 98;
razn_h_mem[7244] = 228;
razn_h_mem[7245] = 104;
razn_h_mem[7246] = 234;
razn_h_mem[7247] = 110;
razn_h_mem[7248] = 240;
razn_h_mem[7249] = 116;
razn_h_mem[7250] = 246;
razn_h_mem[7251] = 122;
razn_h_mem[7252] = 252;
razn_h_mem[7253] = 128;
razn_h_mem[7254] = 4;
razn_h_mem[7255] = 134;
razn_h_mem[7256] = 10;
razn_h_mem[7257] = 140;
razn_h_mem[7258] = 16;
razn_h_mem[7259] = 146;
razn_h_mem[7260] = 22;
razn_h_mem[7261] = 152;
razn_h_mem[7262] = 28;
razn_h_mem[7263] = 158;
razn_h_mem[7264] = 34;
razn_h_mem[7265] = 164;
razn_h_mem[7266] = 40;
razn_h_mem[7267] = 170;
razn_h_mem[7268] = 46;
razn_h_mem[7269] = 176;
razn_h_mem[7270] = 52;
razn_h_mem[7271] = 182;
razn_h_mem[7272] = 58;
razn_h_mem[7273] = 188;
razn_h_mem[7274] = 64;
razn_h_mem[7275] = 194;
razn_h_mem[7276] = 70;
razn_h_mem[7277] = 200;
razn_h_mem[7278] = 76;
razn_h_mem[7279] = 206;
razn_h_mem[7280] = 82;
razn_h_mem[7281] = 212;
razn_h_mem[7282] = 88;
razn_h_mem[7283] = 218;
razn_h_mem[7284] = 94;
razn_h_mem[7285] = 224;
razn_h_mem[7286] = 100;
razn_h_mem[7287] = 230;
razn_h_mem[7288] = 106;
razn_h_mem[7289] = 236;
razn_h_mem[7290] = 112;
razn_h_mem[7291] = 242;
razn_h_mem[7292] = 118;
razn_h_mem[7293] = 248;
razn_h_mem[7294] = 124;
razn_h_mem[7295] = 255;
razn_h_mem[7296] = 0;
razn_h_mem[7297] = 130;
razn_h_mem[7298] = 6;
razn_h_mem[7299] = 136;
razn_h_mem[7300] = 12;
razn_h_mem[7301] = 142;
razn_h_mem[7302] = 18;
razn_h_mem[7303] = 148;
razn_h_mem[7304] = 24;
razn_h_mem[7305] = 154;
razn_h_mem[7306] = 30;
razn_h_mem[7307] = 160;
razn_h_mem[7308] = 36;
razn_h_mem[7309] = 166;
razn_h_mem[7310] = 42;
razn_h_mem[7311] = 172;
razn_h_mem[7312] = 48;
razn_h_mem[7313] = 178;
razn_h_mem[7314] = 54;
razn_h_mem[7315] = 184;
razn_h_mem[7316] = 60;
razn_h_mem[7317] = 190;
razn_h_mem[7318] = 66;
razn_h_mem[7319] = 196;
razn_h_mem[7320] = 72;
razn_h_mem[7321] = 202;
razn_h_mem[7322] = 78;
razn_h_mem[7323] = 208;
razn_h_mem[7324] = 84;
razn_h_mem[7325] = 214;
razn_h_mem[7326] = 90;
razn_h_mem[7327] = 220;
razn_h_mem[7328] = 96;
razn_h_mem[7329] = 226;
razn_h_mem[7330] = 102;
razn_h_mem[7331] = 232;
razn_h_mem[7332] = 108;
razn_h_mem[7333] = 238;
razn_h_mem[7334] = 114;
razn_h_mem[7335] = 244;
razn_h_mem[7336] = 120;
razn_h_mem[7337] = 250;
razn_h_mem[7338] = 126;
razn_h_mem[7339] = 2;
razn_h_mem[7340] = 132;
razn_h_mem[7341] = 8;
razn_h_mem[7342] = 138;
razn_h_mem[7343] = 14;
razn_h_mem[7344] = 144;
razn_h_mem[7345] = 20;
razn_h_mem[7346] = 150;
razn_h_mem[7347] = 26;
razn_h_mem[7348] = 156;
razn_h_mem[7349] = 32;
razn_h_mem[7350] = 162;
razn_h_mem[7351] = 38;
razn_h_mem[7352] = 168;
razn_h_mem[7353] = 44;
razn_h_mem[7354] = 174;
razn_h_mem[7355] = 50;
razn_h_mem[7356] = 180;
razn_h_mem[7357] = 56;
razn_h_mem[7358] = 186;
razn_h_mem[7359] = 62;
razn_h_mem[7360] = 192;
razn_h_mem[7361] = 68;
razn_h_mem[7362] = 198;
razn_h_mem[7363] = 74;
razn_h_mem[7364] = 204;
razn_h_mem[7365] = 80;
razn_h_mem[7366] = 210;
razn_h_mem[7367] = 86;
razn_h_mem[7368] = 216;
razn_h_mem[7369] = 92;
razn_h_mem[7370] = 222;
razn_h_mem[7371] = 98;
razn_h_mem[7372] = 228;
razn_h_mem[7373] = 104;
razn_h_mem[7374] = 234;
razn_h_mem[7375] = 110;
razn_h_mem[7376] = 240;
razn_h_mem[7377] = 116;
razn_h_mem[7378] = 246;
razn_h_mem[7379] = 122;
razn_h_mem[7380] = 252;
razn_h_mem[7381] = 128;
razn_h_mem[7382] = 4;
razn_h_mem[7383] = 134;
razn_h_mem[7384] = 10;
razn_h_mem[7385] = 140;
razn_h_mem[7386] = 16;
razn_h_mem[7387] = 146;
razn_h_mem[7388] = 22;
razn_h_mem[7389] = 152;
razn_h_mem[7390] = 28;
razn_h_mem[7391] = 158;
razn_h_mem[7392] = 34;
razn_h_mem[7393] = 164;
razn_h_mem[7394] = 40;
razn_h_mem[7395] = 170;
razn_h_mem[7396] = 46;
razn_h_mem[7397] = 176;
razn_h_mem[7398] = 52;
razn_h_mem[7399] = 182;
razn_h_mem[7400] = 58;
razn_h_mem[7401] = 188;
razn_h_mem[7402] = 64;
razn_h_mem[7403] = 194;
razn_h_mem[7404] = 70;
razn_h_mem[7405] = 200;
razn_h_mem[7406] = 76;
razn_h_mem[7407] = 206;
razn_h_mem[7408] = 82;
razn_h_mem[7409] = 212;
razn_h_mem[7410] = 88;
razn_h_mem[7411] = 218;
razn_h_mem[7412] = 94;
razn_h_mem[7413] = 224;
razn_h_mem[7414] = 100;
razn_h_mem[7415] = 230;
razn_h_mem[7416] = 106;
razn_h_mem[7417] = 236;
razn_h_mem[7418] = 112;
razn_h_mem[7419] = 242;
razn_h_mem[7420] = 118;
razn_h_mem[7421] = 248;
razn_h_mem[7422] = 124;
razn_h_mem[7423] = 255;
razn_h_mem[7424] = 0;
razn_h_mem[7425] = 130;
razn_h_mem[7426] = 6;
razn_h_mem[7427] = 136;
razn_h_mem[7428] = 12;
razn_h_mem[7429] = 142;
razn_h_mem[7430] = 18;
razn_h_mem[7431] = 148;
razn_h_mem[7432] = 24;
razn_h_mem[7433] = 154;
razn_h_mem[7434] = 30;
razn_h_mem[7435] = 160;
razn_h_mem[7436] = 36;
razn_h_mem[7437] = 166;
razn_h_mem[7438] = 42;
razn_h_mem[7439] = 172;
razn_h_mem[7440] = 48;
razn_h_mem[7441] = 178;
razn_h_mem[7442] = 54;
razn_h_mem[7443] = 184;
razn_h_mem[7444] = 60;
razn_h_mem[7445] = 190;
razn_h_mem[7446] = 66;
razn_h_mem[7447] = 196;
razn_h_mem[7448] = 72;
razn_h_mem[7449] = 202;
razn_h_mem[7450] = 78;
razn_h_mem[7451] = 208;
razn_h_mem[7452] = 84;
razn_h_mem[7453] = 214;
razn_h_mem[7454] = 90;
razn_h_mem[7455] = 220;
razn_h_mem[7456] = 96;
razn_h_mem[7457] = 226;
razn_h_mem[7458] = 102;
razn_h_mem[7459] = 232;
razn_h_mem[7460] = 108;
razn_h_mem[7461] = 238;
razn_h_mem[7462] = 114;
razn_h_mem[7463] = 244;
razn_h_mem[7464] = 120;
razn_h_mem[7465] = 250;
razn_h_mem[7466] = 126;
razn_h_mem[7467] = 2;
razn_h_mem[7468] = 132;
razn_h_mem[7469] = 8;
razn_h_mem[7470] = 138;
razn_h_mem[7471] = 14;
razn_h_mem[7472] = 144;
razn_h_mem[7473] = 20;
razn_h_mem[7474] = 150;
razn_h_mem[7475] = 26;
razn_h_mem[7476] = 156;
razn_h_mem[7477] = 32;
razn_h_mem[7478] = 162;
razn_h_mem[7479] = 38;
razn_h_mem[7480] = 168;
razn_h_mem[7481] = 44;
razn_h_mem[7482] = 174;
razn_h_mem[7483] = 50;
razn_h_mem[7484] = 180;
razn_h_mem[7485] = 56;
razn_h_mem[7486] = 186;
razn_h_mem[7487] = 62;
razn_h_mem[7488] = 192;
razn_h_mem[7489] = 68;
razn_h_mem[7490] = 198;
razn_h_mem[7491] = 74;
razn_h_mem[7492] = 204;
razn_h_mem[7493] = 80;
razn_h_mem[7494] = 210;
razn_h_mem[7495] = 86;
razn_h_mem[7496] = 216;
razn_h_mem[7497] = 92;
razn_h_mem[7498] = 222;
razn_h_mem[7499] = 98;
razn_h_mem[7500] = 228;
razn_h_mem[7501] = 104;
razn_h_mem[7502] = 234;
razn_h_mem[7503] = 110;
razn_h_mem[7504] = 240;
razn_h_mem[7505] = 116;
razn_h_mem[7506] = 246;
razn_h_mem[7507] = 122;
razn_h_mem[7508] = 252;
razn_h_mem[7509] = 128;
razn_h_mem[7510] = 4;
razn_h_mem[7511] = 134;
razn_h_mem[7512] = 10;
razn_h_mem[7513] = 140;
razn_h_mem[7514] = 16;
razn_h_mem[7515] = 146;
razn_h_mem[7516] = 22;
razn_h_mem[7517] = 152;
razn_h_mem[7518] = 28;
razn_h_mem[7519] = 158;
razn_h_mem[7520] = 34;
razn_h_mem[7521] = 164;
razn_h_mem[7522] = 40;
razn_h_mem[7523] = 170;
razn_h_mem[7524] = 46;
razn_h_mem[7525] = 176;
razn_h_mem[7526] = 52;
razn_h_mem[7527] = 182;
razn_h_mem[7528] = 58;
razn_h_mem[7529] = 188;
razn_h_mem[7530] = 64;
razn_h_mem[7531] = 194;
razn_h_mem[7532] = 70;
razn_h_mem[7533] = 200;
razn_h_mem[7534] = 76;
razn_h_mem[7535] = 206;
razn_h_mem[7536] = 82;
razn_h_mem[7537] = 212;
razn_h_mem[7538] = 88;
razn_h_mem[7539] = 218;
razn_h_mem[7540] = 94;
razn_h_mem[7541] = 224;
razn_h_mem[7542] = 100;
razn_h_mem[7543] = 230;
razn_h_mem[7544] = 106;
razn_h_mem[7545] = 236;
razn_h_mem[7546] = 112;
razn_h_mem[7547] = 242;
razn_h_mem[7548] = 118;
razn_h_mem[7549] = 248;
razn_h_mem[7550] = 124;
razn_h_mem[7551] = 255;
razn_h_mem[7552] = 0;
razn_h_mem[7553] = 130;
razn_h_mem[7554] = 6;
razn_h_mem[7555] = 136;
razn_h_mem[7556] = 12;
razn_h_mem[7557] = 142;
razn_h_mem[7558] = 18;
razn_h_mem[7559] = 148;
razn_h_mem[7560] = 24;
razn_h_mem[7561] = 154;
razn_h_mem[7562] = 30;
razn_h_mem[7563] = 160;
razn_h_mem[7564] = 36;
razn_h_mem[7565] = 166;
razn_h_mem[7566] = 42;
razn_h_mem[7567] = 172;
razn_h_mem[7568] = 48;
razn_h_mem[7569] = 178;
razn_h_mem[7570] = 54;
razn_h_mem[7571] = 184;
razn_h_mem[7572] = 60;
razn_h_mem[7573] = 190;
razn_h_mem[7574] = 66;
razn_h_mem[7575] = 196;
razn_h_mem[7576] = 72;
razn_h_mem[7577] = 202;
razn_h_mem[7578] = 78;
razn_h_mem[7579] = 208;
razn_h_mem[7580] = 84;
razn_h_mem[7581] = 214;
razn_h_mem[7582] = 90;
razn_h_mem[7583] = 220;
razn_h_mem[7584] = 96;
razn_h_mem[7585] = 226;
razn_h_mem[7586] = 102;
razn_h_mem[7587] = 232;
razn_h_mem[7588] = 108;
razn_h_mem[7589] = 238;
razn_h_mem[7590] = 114;
razn_h_mem[7591] = 244;
razn_h_mem[7592] = 120;
razn_h_mem[7593] = 250;
razn_h_mem[7594] = 126;
razn_h_mem[7595] = 2;
razn_h_mem[7596] = 132;
razn_h_mem[7597] = 8;
razn_h_mem[7598] = 138;
razn_h_mem[7599] = 14;
razn_h_mem[7600] = 144;
razn_h_mem[7601] = 20;
razn_h_mem[7602] = 150;
razn_h_mem[7603] = 26;
razn_h_mem[7604] = 156;
razn_h_mem[7605] = 32;
razn_h_mem[7606] = 162;
razn_h_mem[7607] = 38;
razn_h_mem[7608] = 168;
razn_h_mem[7609] = 44;
razn_h_mem[7610] = 174;
razn_h_mem[7611] = 50;
razn_h_mem[7612] = 180;
razn_h_mem[7613] = 56;
razn_h_mem[7614] = 186;
razn_h_mem[7615] = 62;
razn_h_mem[7616] = 192;
razn_h_mem[7617] = 68;
razn_h_mem[7618] = 198;
razn_h_mem[7619] = 74;
razn_h_mem[7620] = 204;
razn_h_mem[7621] = 80;
razn_h_mem[7622] = 210;
razn_h_mem[7623] = 86;
razn_h_mem[7624] = 216;
razn_h_mem[7625] = 92;
razn_h_mem[7626] = 222;
razn_h_mem[7627] = 98;
razn_h_mem[7628] = 228;
razn_h_mem[7629] = 104;
razn_h_mem[7630] = 234;
razn_h_mem[7631] = 110;
razn_h_mem[7632] = 240;
razn_h_mem[7633] = 116;
razn_h_mem[7634] = 246;
razn_h_mem[7635] = 122;
razn_h_mem[7636] = 252;
razn_h_mem[7637] = 128;
razn_h_mem[7638] = 4;
razn_h_mem[7639] = 134;
razn_h_mem[7640] = 10;
razn_h_mem[7641] = 140;
razn_h_mem[7642] = 16;
razn_h_mem[7643] = 146;
razn_h_mem[7644] = 22;
razn_h_mem[7645] = 152;
razn_h_mem[7646] = 28;
razn_h_mem[7647] = 158;
razn_h_mem[7648] = 34;
razn_h_mem[7649] = 164;
razn_h_mem[7650] = 40;
razn_h_mem[7651] = 170;
razn_h_mem[7652] = 46;
razn_h_mem[7653] = 176;
razn_h_mem[7654] = 52;
razn_h_mem[7655] = 182;
razn_h_mem[7656] = 58;
razn_h_mem[7657] = 188;
razn_h_mem[7658] = 64;
razn_h_mem[7659] = 194;
razn_h_mem[7660] = 70;
razn_h_mem[7661] = 200;
razn_h_mem[7662] = 76;
razn_h_mem[7663] = 206;
razn_h_mem[7664] = 82;
razn_h_mem[7665] = 212;
razn_h_mem[7666] = 88;
razn_h_mem[7667] = 218;
razn_h_mem[7668] = 94;
razn_h_mem[7669] = 224;
razn_h_mem[7670] = 100;
razn_h_mem[7671] = 230;
razn_h_mem[7672] = 106;
razn_h_mem[7673] = 236;
razn_h_mem[7674] = 112;
razn_h_mem[7675] = 242;
razn_h_mem[7676] = 118;
razn_h_mem[7677] = 248;
razn_h_mem[7678] = 124;
razn_h_mem[7679] = 255;
razn_h_mem[7680] = 0;
razn_h_mem[7681] = 130;
razn_h_mem[7682] = 6;
razn_h_mem[7683] = 136;
razn_h_mem[7684] = 12;
razn_h_mem[7685] = 142;
razn_h_mem[7686] = 18;
razn_h_mem[7687] = 148;
razn_h_mem[7688] = 24;
razn_h_mem[7689] = 154;
razn_h_mem[7690] = 30;
razn_h_mem[7691] = 160;
razn_h_mem[7692] = 36;
razn_h_mem[7693] = 166;
razn_h_mem[7694] = 42;
razn_h_mem[7695] = 172;
razn_h_mem[7696] = 48;
razn_h_mem[7697] = 178;
razn_h_mem[7698] = 54;
razn_h_mem[7699] = 184;
razn_h_mem[7700] = 60;
razn_h_mem[7701] = 190;
razn_h_mem[7702] = 66;
razn_h_mem[7703] = 196;
razn_h_mem[7704] = 72;
razn_h_mem[7705] = 202;
razn_h_mem[7706] = 78;
razn_h_mem[7707] = 208;
razn_h_mem[7708] = 84;
razn_h_mem[7709] = 214;
razn_h_mem[7710] = 90;
razn_h_mem[7711] = 220;
razn_h_mem[7712] = 96;
razn_h_mem[7713] = 226;
razn_h_mem[7714] = 102;
razn_h_mem[7715] = 232;
razn_h_mem[7716] = 108;
razn_h_mem[7717] = 238;
razn_h_mem[7718] = 114;
razn_h_mem[7719] = 244;
razn_h_mem[7720] = 120;
razn_h_mem[7721] = 250;
razn_h_mem[7722] = 126;
razn_h_mem[7723] = 2;
razn_h_mem[7724] = 132;
razn_h_mem[7725] = 8;
razn_h_mem[7726] = 138;
razn_h_mem[7727] = 14;
razn_h_mem[7728] = 144;
razn_h_mem[7729] = 20;
razn_h_mem[7730] = 150;
razn_h_mem[7731] = 26;
razn_h_mem[7732] = 156;
razn_h_mem[7733] = 32;
razn_h_mem[7734] = 162;
razn_h_mem[7735] = 38;
razn_h_mem[7736] = 168;
razn_h_mem[7737] = 44;
razn_h_mem[7738] = 174;
razn_h_mem[7739] = 50;
razn_h_mem[7740] = 180;
razn_h_mem[7741] = 56;
razn_h_mem[7742] = 186;
razn_h_mem[7743] = 62;
razn_h_mem[7744] = 192;
razn_h_mem[7745] = 68;
razn_h_mem[7746] = 198;
razn_h_mem[7747] = 74;
razn_h_mem[7748] = 204;
razn_h_mem[7749] = 80;
razn_h_mem[7750] = 210;
razn_h_mem[7751] = 86;
razn_h_mem[7752] = 216;
razn_h_mem[7753] = 92;
razn_h_mem[7754] = 222;
razn_h_mem[7755] = 98;
razn_h_mem[7756] = 228;
razn_h_mem[7757] = 104;
razn_h_mem[7758] = 234;
razn_h_mem[7759] = 110;
razn_h_mem[7760] = 240;
razn_h_mem[7761] = 116;
razn_h_mem[7762] = 246;
razn_h_mem[7763] = 122;
razn_h_mem[7764] = 252;
razn_h_mem[7765] = 128;
razn_h_mem[7766] = 4;
razn_h_mem[7767] = 134;
razn_h_mem[7768] = 10;
razn_h_mem[7769] = 140;
razn_h_mem[7770] = 16;
razn_h_mem[7771] = 146;
razn_h_mem[7772] = 22;
razn_h_mem[7773] = 152;
razn_h_mem[7774] = 28;
razn_h_mem[7775] = 158;
razn_h_mem[7776] = 34;
razn_h_mem[7777] = 164;
razn_h_mem[7778] = 40;
razn_h_mem[7779] = 170;
razn_h_mem[7780] = 46;
razn_h_mem[7781] = 176;
razn_h_mem[7782] = 52;
razn_h_mem[7783] = 182;
razn_h_mem[7784] = 58;
razn_h_mem[7785] = 188;
razn_h_mem[7786] = 64;
razn_h_mem[7787] = 194;
razn_h_mem[7788] = 70;
razn_h_mem[7789] = 200;
razn_h_mem[7790] = 76;
razn_h_mem[7791] = 206;
razn_h_mem[7792] = 82;
razn_h_mem[7793] = 212;
razn_h_mem[7794] = 88;
razn_h_mem[7795] = 218;
razn_h_mem[7796] = 94;
razn_h_mem[7797] = 224;
razn_h_mem[7798] = 100;
razn_h_mem[7799] = 230;
razn_h_mem[7800] = 106;
razn_h_mem[7801] = 236;
razn_h_mem[7802] = 112;
razn_h_mem[7803] = 242;
razn_h_mem[7804] = 118;
razn_h_mem[7805] = 248;
razn_h_mem[7806] = 124;
razn_h_mem[7807] = 255;
razn_h_mem[7808] = 0;
razn_h_mem[7809] = 130;
razn_h_mem[7810] = 6;
razn_h_mem[7811] = 136;
razn_h_mem[7812] = 12;
razn_h_mem[7813] = 142;
razn_h_mem[7814] = 18;
razn_h_mem[7815] = 148;
razn_h_mem[7816] = 24;
razn_h_mem[7817] = 154;
razn_h_mem[7818] = 30;
razn_h_mem[7819] = 160;
razn_h_mem[7820] = 36;
razn_h_mem[7821] = 166;
razn_h_mem[7822] = 42;
razn_h_mem[7823] = 172;
razn_h_mem[7824] = 48;
razn_h_mem[7825] = 178;
razn_h_mem[7826] = 54;
razn_h_mem[7827] = 184;
razn_h_mem[7828] = 60;
razn_h_mem[7829] = 190;
razn_h_mem[7830] = 66;
razn_h_mem[7831] = 196;
razn_h_mem[7832] = 72;
razn_h_mem[7833] = 202;
razn_h_mem[7834] = 78;
razn_h_mem[7835] = 208;
razn_h_mem[7836] = 84;
razn_h_mem[7837] = 214;
razn_h_mem[7838] = 90;
razn_h_mem[7839] = 220;
razn_h_mem[7840] = 96;
razn_h_mem[7841] = 226;
razn_h_mem[7842] = 102;
razn_h_mem[7843] = 232;
razn_h_mem[7844] = 108;
razn_h_mem[7845] = 238;
razn_h_mem[7846] = 114;
razn_h_mem[7847] = 244;
razn_h_mem[7848] = 120;
razn_h_mem[7849] = 250;
razn_h_mem[7850] = 126;
razn_h_mem[7851] = 2;
razn_h_mem[7852] = 132;
razn_h_mem[7853] = 8;
razn_h_mem[7854] = 138;
razn_h_mem[7855] = 14;
razn_h_mem[7856] = 144;
razn_h_mem[7857] = 20;
razn_h_mem[7858] = 150;
razn_h_mem[7859] = 26;
razn_h_mem[7860] = 156;
razn_h_mem[7861] = 32;
razn_h_mem[7862] = 162;
razn_h_mem[7863] = 38;
razn_h_mem[7864] = 168;
razn_h_mem[7865] = 44;
razn_h_mem[7866] = 174;
razn_h_mem[7867] = 50;
razn_h_mem[7868] = 180;
razn_h_mem[7869] = 56;
razn_h_mem[7870] = 186;
razn_h_mem[7871] = 62;
razn_h_mem[7872] = 192;
razn_h_mem[7873] = 68;
razn_h_mem[7874] = 198;
razn_h_mem[7875] = 74;
razn_h_mem[7876] = 204;
razn_h_mem[7877] = 80;
razn_h_mem[7878] = 210;
razn_h_mem[7879] = 86;
razn_h_mem[7880] = 216;
razn_h_mem[7881] = 92;
razn_h_mem[7882] = 222;
razn_h_mem[7883] = 98;
razn_h_mem[7884] = 228;
razn_h_mem[7885] = 104;
razn_h_mem[7886] = 234;
razn_h_mem[7887] = 110;
razn_h_mem[7888] = 240;
razn_h_mem[7889] = 116;
razn_h_mem[7890] = 246;
razn_h_mem[7891] = 122;
razn_h_mem[7892] = 252;
razn_h_mem[7893] = 128;
razn_h_mem[7894] = 4;
razn_h_mem[7895] = 134;
razn_h_mem[7896] = 10;
razn_h_mem[7897] = 140;
razn_h_mem[7898] = 16;
razn_h_mem[7899] = 146;
razn_h_mem[7900] = 22;
razn_h_mem[7901] = 152;
razn_h_mem[7902] = 28;
razn_h_mem[7903] = 158;
razn_h_mem[7904] = 34;
razn_h_mem[7905] = 164;
razn_h_mem[7906] = 40;
razn_h_mem[7907] = 170;
razn_h_mem[7908] = 46;
razn_h_mem[7909] = 176;
razn_h_mem[7910] = 52;
razn_h_mem[7911] = 182;
razn_h_mem[7912] = 58;
razn_h_mem[7913] = 188;
razn_h_mem[7914] = 64;
razn_h_mem[7915] = 194;
razn_h_mem[7916] = 70;
razn_h_mem[7917] = 200;
razn_h_mem[7918] = 76;
razn_h_mem[7919] = 206;
razn_h_mem[7920] = 82;
razn_h_mem[7921] = 212;
razn_h_mem[7922] = 88;
razn_h_mem[7923] = 218;
razn_h_mem[7924] = 94;
razn_h_mem[7925] = 224;
razn_h_mem[7926] = 100;
razn_h_mem[7927] = 230;
razn_h_mem[7928] = 106;
razn_h_mem[7929] = 236;
razn_h_mem[7930] = 112;
razn_h_mem[7931] = 242;
razn_h_mem[7932] = 118;
razn_h_mem[7933] = 248;
razn_h_mem[7934] = 124;
razn_h_mem[7935] = 255;
razn_h_mem[7936] = 0;
razn_h_mem[7937] = 130;
razn_h_mem[7938] = 6;
razn_h_mem[7939] = 136;
razn_h_mem[7940] = 12;
razn_h_mem[7941] = 142;
razn_h_mem[7942] = 18;
razn_h_mem[7943] = 148;
razn_h_mem[7944] = 24;
razn_h_mem[7945] = 154;
razn_h_mem[7946] = 30;
razn_h_mem[7947] = 160;
razn_h_mem[7948] = 36;
razn_h_mem[7949] = 166;
razn_h_mem[7950] = 42;
razn_h_mem[7951] = 172;
razn_h_mem[7952] = 48;
razn_h_mem[7953] = 178;
razn_h_mem[7954] = 54;
razn_h_mem[7955] = 184;
razn_h_mem[7956] = 60;
razn_h_mem[7957] = 190;
razn_h_mem[7958] = 66;
razn_h_mem[7959] = 196;
razn_h_mem[7960] = 72;
razn_h_mem[7961] = 202;
razn_h_mem[7962] = 78;
razn_h_mem[7963] = 208;
razn_h_mem[7964] = 84;
razn_h_mem[7965] = 214;
razn_h_mem[7966] = 90;
razn_h_mem[7967] = 220;
razn_h_mem[7968] = 96;
razn_h_mem[7969] = 226;
razn_h_mem[7970] = 102;
razn_h_mem[7971] = 232;
razn_h_mem[7972] = 108;
razn_h_mem[7973] = 238;
razn_h_mem[7974] = 114;
razn_h_mem[7975] = 244;
razn_h_mem[7976] = 120;
razn_h_mem[7977] = 250;
razn_h_mem[7978] = 126;
razn_h_mem[7979] = 2;
razn_h_mem[7980] = 132;
razn_h_mem[7981] = 8;
razn_h_mem[7982] = 138;
razn_h_mem[7983] = 14;
razn_h_mem[7984] = 144;
razn_h_mem[7985] = 20;
razn_h_mem[7986] = 150;
razn_h_mem[7987] = 26;
razn_h_mem[7988] = 156;
razn_h_mem[7989] = 32;
razn_h_mem[7990] = 162;
razn_h_mem[7991] = 38;
razn_h_mem[7992] = 168;
razn_h_mem[7993] = 44;
razn_h_mem[7994] = 174;
razn_h_mem[7995] = 50;
razn_h_mem[7996] = 180;
razn_h_mem[7997] = 56;
razn_h_mem[7998] = 186;
razn_h_mem[7999] = 62;
razn_h_mem[8000] = 192;
razn_h_mem[8001] = 68;
razn_h_mem[8002] = 198;
razn_h_mem[8003] = 74;
razn_h_mem[8004] = 204;
razn_h_mem[8005] = 80;
razn_h_mem[8006] = 210;
razn_h_mem[8007] = 86;
razn_h_mem[8008] = 216;
razn_h_mem[8009] = 92;
razn_h_mem[8010] = 222;
razn_h_mem[8011] = 98;
razn_h_mem[8012] = 228;
razn_h_mem[8013] = 104;
razn_h_mem[8014] = 234;
razn_h_mem[8015] = 110;
razn_h_mem[8016] = 240;
razn_h_mem[8017] = 116;
razn_h_mem[8018] = 246;
razn_h_mem[8019] = 122;
razn_h_mem[8020] = 252;
razn_h_mem[8021] = 128;
razn_h_mem[8022] = 4;
razn_h_mem[8023] = 134;
razn_h_mem[8024] = 10;
razn_h_mem[8025] = 140;
razn_h_mem[8026] = 16;
razn_h_mem[8027] = 146;
razn_h_mem[8028] = 22;
razn_h_mem[8029] = 152;
razn_h_mem[8030] = 28;
razn_h_mem[8031] = 158;
razn_h_mem[8032] = 34;
razn_h_mem[8033] = 164;
razn_h_mem[8034] = 40;
razn_h_mem[8035] = 170;
razn_h_mem[8036] = 46;
razn_h_mem[8037] = 176;
razn_h_mem[8038] = 52;
razn_h_mem[8039] = 182;
razn_h_mem[8040] = 58;
razn_h_mem[8041] = 188;
razn_h_mem[8042] = 64;
razn_h_mem[8043] = 194;
razn_h_mem[8044] = 70;
razn_h_mem[8045] = 200;
razn_h_mem[8046] = 76;
razn_h_mem[8047] = 206;
razn_h_mem[8048] = 82;
razn_h_mem[8049] = 212;
razn_h_mem[8050] = 88;
razn_h_mem[8051] = 218;
razn_h_mem[8052] = 94;
razn_h_mem[8053] = 224;
razn_h_mem[8054] = 100;
razn_h_mem[8055] = 230;
razn_h_mem[8056] = 106;
razn_h_mem[8057] = 236;
razn_h_mem[8058] = 112;
razn_h_mem[8059] = 242;
razn_h_mem[8060] = 118;
razn_h_mem[8061] = 248;
razn_h_mem[8062] = 124;
razn_h_mem[8063] = 255;
razn_h_mem[8064] = 0;
razn_h_mem[8065] = 130;
razn_h_mem[8066] = 6;
razn_h_mem[8067] = 136;
razn_h_mem[8068] = 12;
razn_h_mem[8069] = 142;
razn_h_mem[8070] = 18;
razn_h_mem[8071] = 148;
razn_h_mem[8072] = 24;
razn_h_mem[8073] = 154;
razn_h_mem[8074] = 30;
razn_h_mem[8075] = 160;
razn_h_mem[8076] = 36;
razn_h_mem[8077] = 166;
razn_h_mem[8078] = 42;
razn_h_mem[8079] = 172;
razn_h_mem[8080] = 48;
razn_h_mem[8081] = 178;
razn_h_mem[8082] = 54;
razn_h_mem[8083] = 184;
razn_h_mem[8084] = 60;
razn_h_mem[8085] = 190;
razn_h_mem[8086] = 66;
razn_h_mem[8087] = 196;
razn_h_mem[8088] = 72;
razn_h_mem[8089] = 202;
razn_h_mem[8090] = 78;
razn_h_mem[8091] = 208;
razn_h_mem[8092] = 84;
razn_h_mem[8093] = 214;
razn_h_mem[8094] = 90;
razn_h_mem[8095] = 220;
razn_h_mem[8096] = 96;
razn_h_mem[8097] = 226;
razn_h_mem[8098] = 102;
razn_h_mem[8099] = 232;
razn_h_mem[8100] = 108;
razn_h_mem[8101] = 238;
razn_h_mem[8102] = 114;
razn_h_mem[8103] = 244;
razn_h_mem[8104] = 120;
razn_h_mem[8105] = 250;
razn_h_mem[8106] = 126;
razn_h_mem[8107] = 2;
razn_h_mem[8108] = 132;
razn_h_mem[8109] = 8;
razn_h_mem[8110] = 138;
razn_h_mem[8111] = 14;
razn_h_mem[8112] = 144;
razn_h_mem[8113] = 20;
razn_h_mem[8114] = 150;
razn_h_mem[8115] = 26;
razn_h_mem[8116] = 156;
razn_h_mem[8117] = 32;
razn_h_mem[8118] = 162;
razn_h_mem[8119] = 38;
razn_h_mem[8120] = 168;
razn_h_mem[8121] = 44;
razn_h_mem[8122] = 174;
razn_h_mem[8123] = 50;
razn_h_mem[8124] = 180;
razn_h_mem[8125] = 56;
razn_h_mem[8126] = 186;
razn_h_mem[8127] = 62;
razn_h_mem[8128] = 192;
razn_h_mem[8129] = 68;
razn_h_mem[8130] = 198;
razn_h_mem[8131] = 74;
razn_h_mem[8132] = 204;
razn_h_mem[8133] = 80;
razn_h_mem[8134] = 210;
razn_h_mem[8135] = 86;
razn_h_mem[8136] = 216;
razn_h_mem[8137] = 92;
razn_h_mem[8138] = 222;
razn_h_mem[8139] = 98;
razn_h_mem[8140] = 228;
razn_h_mem[8141] = 104;
razn_h_mem[8142] = 234;
razn_h_mem[8143] = 110;
razn_h_mem[8144] = 240;
razn_h_mem[8145] = 116;
razn_h_mem[8146] = 246;
razn_h_mem[8147] = 122;
razn_h_mem[8148] = 252;
razn_h_mem[8149] = 128;
razn_h_mem[8150] = 4;
razn_h_mem[8151] = 134;
razn_h_mem[8152] = 10;
razn_h_mem[8153] = 140;
razn_h_mem[8154] = 16;
razn_h_mem[8155] = 146;
razn_h_mem[8156] = 22;
razn_h_mem[8157] = 152;
razn_h_mem[8158] = 28;
razn_h_mem[8159] = 158;
razn_h_mem[8160] = 34;
razn_h_mem[8161] = 164;
razn_h_mem[8162] = 40;
razn_h_mem[8163] = 170;
razn_h_mem[8164] = 46;
razn_h_mem[8165] = 176;
razn_h_mem[8166] = 52;
razn_h_mem[8167] = 182;
razn_h_mem[8168] = 58;
razn_h_mem[8169] = 188;
razn_h_mem[8170] = 64;
razn_h_mem[8171] = 194;
razn_h_mem[8172] = 70;
razn_h_mem[8173] = 200;
razn_h_mem[8174] = 76;
razn_h_mem[8175] = 206;
razn_h_mem[8176] = 82;
razn_h_mem[8177] = 212;
razn_h_mem[8178] = 88;
razn_h_mem[8179] = 218;
razn_h_mem[8180] = 94;
razn_h_mem[8181] = 224;
razn_h_mem[8182] = 100;
razn_h_mem[8183] = 230;
razn_h_mem[8184] = 106;
razn_h_mem[8185] = 236;
razn_h_mem[8186] = 112;
razn_h_mem[8187] = 242;
razn_h_mem[8188] = 118;
razn_h_mem[8189] = 248;
razn_h_mem[8190] = 124;
razn_h_mem[8191] = 255;
razn_h_mem[8192] = 0;
razn_h_mem[8193] = 130;
razn_h_mem[8194] = 6;
razn_h_mem[8195] = 136;
razn_h_mem[8196] = 12;
razn_h_mem[8197] = 142;
razn_h_mem[8198] = 18;
razn_h_mem[8199] = 148;
razn_h_mem[8200] = 24;
razn_h_mem[8201] = 154;
razn_h_mem[8202] = 30;
razn_h_mem[8203] = 160;
razn_h_mem[8204] = 36;
razn_h_mem[8205] = 166;
razn_h_mem[8206] = 42;
razn_h_mem[8207] = 172;
razn_h_mem[8208] = 48;
razn_h_mem[8209] = 178;
razn_h_mem[8210] = 54;
razn_h_mem[8211] = 184;
razn_h_mem[8212] = 60;
razn_h_mem[8213] = 190;
razn_h_mem[8214] = 66;
razn_h_mem[8215] = 196;
razn_h_mem[8216] = 72;
razn_h_mem[8217] = 202;
razn_h_mem[8218] = 78;
razn_h_mem[8219] = 208;
razn_h_mem[8220] = 84;
razn_h_mem[8221] = 214;
razn_h_mem[8222] = 90;
razn_h_mem[8223] = 220;
razn_h_mem[8224] = 96;
razn_h_mem[8225] = 226;
razn_h_mem[8226] = 102;
razn_h_mem[8227] = 232;
razn_h_mem[8228] = 108;
razn_h_mem[8229] = 238;
razn_h_mem[8230] = 114;
razn_h_mem[8231] = 244;
razn_h_mem[8232] = 120;
razn_h_mem[8233] = 250;
razn_h_mem[8234] = 126;
razn_h_mem[8235] = 2;
razn_h_mem[8236] = 132;
razn_h_mem[8237] = 8;
razn_h_mem[8238] = 138;
razn_h_mem[8239] = 14;
razn_h_mem[8240] = 144;
razn_h_mem[8241] = 20;
razn_h_mem[8242] = 150;
razn_h_mem[8243] = 26;
razn_h_mem[8244] = 156;
razn_h_mem[8245] = 32;
razn_h_mem[8246] = 162;
razn_h_mem[8247] = 38;
razn_h_mem[8248] = 168;
razn_h_mem[8249] = 44;
razn_h_mem[8250] = 174;
razn_h_mem[8251] = 50;
razn_h_mem[8252] = 180;
razn_h_mem[8253] = 56;
razn_h_mem[8254] = 186;
razn_h_mem[8255] = 62;
razn_h_mem[8256] = 192;
razn_h_mem[8257] = 68;
razn_h_mem[8258] = 198;
razn_h_mem[8259] = 74;
razn_h_mem[8260] = 204;
razn_h_mem[8261] = 80;
razn_h_mem[8262] = 210;
razn_h_mem[8263] = 86;
razn_h_mem[8264] = 216;
razn_h_mem[8265] = 92;
razn_h_mem[8266] = 222;
razn_h_mem[8267] = 98;
razn_h_mem[8268] = 228;
razn_h_mem[8269] = 104;
razn_h_mem[8270] = 234;
razn_h_mem[8271] = 110;
razn_h_mem[8272] = 240;
razn_h_mem[8273] = 116;
razn_h_mem[8274] = 246;
razn_h_mem[8275] = 122;
razn_h_mem[8276] = 252;
razn_h_mem[8277] = 128;
razn_h_mem[8278] = 4;
razn_h_mem[8279] = 134;
razn_h_mem[8280] = 10;
razn_h_mem[8281] = 140;
razn_h_mem[8282] = 16;
razn_h_mem[8283] = 146;
razn_h_mem[8284] = 22;
razn_h_mem[8285] = 152;
razn_h_mem[8286] = 28;
razn_h_mem[8287] = 158;
razn_h_mem[8288] = 34;
razn_h_mem[8289] = 164;
razn_h_mem[8290] = 40;
razn_h_mem[8291] = 170;
razn_h_mem[8292] = 46;
razn_h_mem[8293] = 176;
razn_h_mem[8294] = 52;
razn_h_mem[8295] = 182;
razn_h_mem[8296] = 58;
razn_h_mem[8297] = 188;
razn_h_mem[8298] = 64;
razn_h_mem[8299] = 194;
razn_h_mem[8300] = 70;
razn_h_mem[8301] = 200;
razn_h_mem[8302] = 76;
razn_h_mem[8303] = 206;
razn_h_mem[8304] = 82;
razn_h_mem[8305] = 212;
razn_h_mem[8306] = 88;
razn_h_mem[8307] = 218;
razn_h_mem[8308] = 94;
razn_h_mem[8309] = 224;
razn_h_mem[8310] = 100;
razn_h_mem[8311] = 230;
razn_h_mem[8312] = 106;
razn_h_mem[8313] = 236;
razn_h_mem[8314] = 112;
razn_h_mem[8315] = 242;
razn_h_mem[8316] = 118;
razn_h_mem[8317] = 248;
razn_h_mem[8318] = 124;
razn_h_mem[8319] = 255;
razn_h_mem[8320] = 0;
razn_h_mem[8321] = 130;
razn_h_mem[8322] = 6;
razn_h_mem[8323] = 136;
razn_h_mem[8324] = 12;
razn_h_mem[8325] = 142;
razn_h_mem[8326] = 18;
razn_h_mem[8327] = 148;
razn_h_mem[8328] = 24;
razn_h_mem[8329] = 154;
razn_h_mem[8330] = 30;
razn_h_mem[8331] = 160;
razn_h_mem[8332] = 36;
razn_h_mem[8333] = 166;
razn_h_mem[8334] = 42;
razn_h_mem[8335] = 172;
razn_h_mem[8336] = 48;
razn_h_mem[8337] = 178;
razn_h_mem[8338] = 54;
razn_h_mem[8339] = 184;
razn_h_mem[8340] = 60;
razn_h_mem[8341] = 190;
razn_h_mem[8342] = 66;
razn_h_mem[8343] = 196;
razn_h_mem[8344] = 72;
razn_h_mem[8345] = 202;
razn_h_mem[8346] = 78;
razn_h_mem[8347] = 208;
razn_h_mem[8348] = 84;
razn_h_mem[8349] = 214;
razn_h_mem[8350] = 90;
razn_h_mem[8351] = 220;
razn_h_mem[8352] = 96;
razn_h_mem[8353] = 226;
razn_h_mem[8354] = 102;
razn_h_mem[8355] = 232;
razn_h_mem[8356] = 108;
razn_h_mem[8357] = 238;
razn_h_mem[8358] = 114;
razn_h_mem[8359] = 244;
razn_h_mem[8360] = 120;
razn_h_mem[8361] = 250;
razn_h_mem[8362] = 126;
razn_h_mem[8363] = 2;
razn_h_mem[8364] = 132;
razn_h_mem[8365] = 8;
razn_h_mem[8366] = 138;
razn_h_mem[8367] = 14;
razn_h_mem[8368] = 144;
razn_h_mem[8369] = 20;
razn_h_mem[8370] = 150;
razn_h_mem[8371] = 26;
razn_h_mem[8372] = 156;
razn_h_mem[8373] = 32;
razn_h_mem[8374] = 162;
razn_h_mem[8375] = 38;
razn_h_mem[8376] = 168;
razn_h_mem[8377] = 44;
razn_h_mem[8378] = 174;
razn_h_mem[8379] = 50;
razn_h_mem[8380] = 180;
razn_h_mem[8381] = 56;
razn_h_mem[8382] = 186;
razn_h_mem[8383] = 62;
razn_h_mem[8384] = 192;
razn_h_mem[8385] = 68;
razn_h_mem[8386] = 198;
razn_h_mem[8387] = 74;
razn_h_mem[8388] = 204;
razn_h_mem[8389] = 80;
razn_h_mem[8390] = 210;
razn_h_mem[8391] = 86;
razn_h_mem[8392] = 216;
razn_h_mem[8393] = 92;
razn_h_mem[8394] = 222;
razn_h_mem[8395] = 98;
razn_h_mem[8396] = 228;
razn_h_mem[8397] = 104;
razn_h_mem[8398] = 234;
razn_h_mem[8399] = 110;
razn_h_mem[8400] = 240;
razn_h_mem[8401] = 116;
razn_h_mem[8402] = 246;
razn_h_mem[8403] = 122;
razn_h_mem[8404] = 252;
razn_h_mem[8405] = 128;
razn_h_mem[8406] = 4;
razn_h_mem[8407] = 134;
razn_h_mem[8408] = 10;
razn_h_mem[8409] = 140;
razn_h_mem[8410] = 16;
razn_h_mem[8411] = 146;
razn_h_mem[8412] = 22;
razn_h_mem[8413] = 152;
razn_h_mem[8414] = 28;
razn_h_mem[8415] = 158;
razn_h_mem[8416] = 34;
razn_h_mem[8417] = 164;
razn_h_mem[8418] = 40;
razn_h_mem[8419] = 170;
razn_h_mem[8420] = 46;
razn_h_mem[8421] = 176;
razn_h_mem[8422] = 52;
razn_h_mem[8423] = 182;
razn_h_mem[8424] = 58;
razn_h_mem[8425] = 188;
razn_h_mem[8426] = 64;
razn_h_mem[8427] = 194;
razn_h_mem[8428] = 70;
razn_h_mem[8429] = 200;
razn_h_mem[8430] = 76;
razn_h_mem[8431] = 206;
razn_h_mem[8432] = 82;
razn_h_mem[8433] = 212;
razn_h_mem[8434] = 88;
razn_h_mem[8435] = 218;
razn_h_mem[8436] = 94;
razn_h_mem[8437] = 224;
razn_h_mem[8438] = 100;
razn_h_mem[8439] = 230;
razn_h_mem[8440] = 106;
razn_h_mem[8441] = 236;
razn_h_mem[8442] = 112;
razn_h_mem[8443] = 242;
razn_h_mem[8444] = 118;
razn_h_mem[8445] = 248;
razn_h_mem[8446] = 124;
razn_h_mem[8447] = 255;
razn_h_mem[8448] = 0;
razn_h_mem[8449] = 130;
razn_h_mem[8450] = 6;
razn_h_mem[8451] = 136;
razn_h_mem[8452] = 12;
razn_h_mem[8453] = 142;
razn_h_mem[8454] = 18;
razn_h_mem[8455] = 148;
razn_h_mem[8456] = 24;
razn_h_mem[8457] = 154;
razn_h_mem[8458] = 30;
razn_h_mem[8459] = 160;
razn_h_mem[8460] = 36;
razn_h_mem[8461] = 166;
razn_h_mem[8462] = 42;
razn_h_mem[8463] = 172;
razn_h_mem[8464] = 48;
razn_h_mem[8465] = 178;
razn_h_mem[8466] = 54;
razn_h_mem[8467] = 184;
razn_h_mem[8468] = 60;
razn_h_mem[8469] = 190;
razn_h_mem[8470] = 66;
razn_h_mem[8471] = 196;
razn_h_mem[8472] = 72;
razn_h_mem[8473] = 202;
razn_h_mem[8474] = 78;
razn_h_mem[8475] = 208;
razn_h_mem[8476] = 84;
razn_h_mem[8477] = 214;
razn_h_mem[8478] = 90;
razn_h_mem[8479] = 220;
razn_h_mem[8480] = 96;
razn_h_mem[8481] = 226;
razn_h_mem[8482] = 102;
razn_h_mem[8483] = 232;
razn_h_mem[8484] = 108;
razn_h_mem[8485] = 238;
razn_h_mem[8486] = 114;
razn_h_mem[8487] = 244;
razn_h_mem[8488] = 120;
razn_h_mem[8489] = 250;
razn_h_mem[8490] = 126;
razn_h_mem[8491] = 2;
razn_h_mem[8492] = 132;
razn_h_mem[8493] = 8;
razn_h_mem[8494] = 138;
razn_h_mem[8495] = 14;
razn_h_mem[8496] = 144;
razn_h_mem[8497] = 20;
razn_h_mem[8498] = 150;
razn_h_mem[8499] = 26;
razn_h_mem[8500] = 156;
razn_h_mem[8501] = 32;
razn_h_mem[8502] = 162;
razn_h_mem[8503] = 38;
razn_h_mem[8504] = 168;
razn_h_mem[8505] = 44;
razn_h_mem[8506] = 174;
razn_h_mem[8507] = 50;
razn_h_mem[8508] = 180;
razn_h_mem[8509] = 56;
razn_h_mem[8510] = 186;
razn_h_mem[8511] = 62;
razn_h_mem[8512] = 192;
razn_h_mem[8513] = 68;
razn_h_mem[8514] = 198;
razn_h_mem[8515] = 74;
razn_h_mem[8516] = 204;
razn_h_mem[8517] = 80;
razn_h_mem[8518] = 210;
razn_h_mem[8519] = 86;
razn_h_mem[8520] = 216;
razn_h_mem[8521] = 92;
razn_h_mem[8522] = 222;
razn_h_mem[8523] = 98;
razn_h_mem[8524] = 228;
razn_h_mem[8525] = 104;
razn_h_mem[8526] = 234;
razn_h_mem[8527] = 110;
razn_h_mem[8528] = 240;
razn_h_mem[8529] = 116;
razn_h_mem[8530] = 246;
razn_h_mem[8531] = 122;
razn_h_mem[8532] = 252;
razn_h_mem[8533] = 128;
razn_h_mem[8534] = 4;
razn_h_mem[8535] = 134;
razn_h_mem[8536] = 10;
razn_h_mem[8537] = 140;
razn_h_mem[8538] = 16;
razn_h_mem[8539] = 146;
razn_h_mem[8540] = 22;
razn_h_mem[8541] = 152;
razn_h_mem[8542] = 28;
razn_h_mem[8543] = 158;
razn_h_mem[8544] = 34;
razn_h_mem[8545] = 164;
razn_h_mem[8546] = 40;
razn_h_mem[8547] = 170;
razn_h_mem[8548] = 46;
razn_h_mem[8549] = 176;
razn_h_mem[8550] = 52;
razn_h_mem[8551] = 182;
razn_h_mem[8552] = 58;
razn_h_mem[8553] = 188;
razn_h_mem[8554] = 64;
razn_h_mem[8555] = 194;
razn_h_mem[8556] = 70;
razn_h_mem[8557] = 200;
razn_h_mem[8558] = 76;
razn_h_mem[8559] = 206;
razn_h_mem[8560] = 82;
razn_h_mem[8561] = 212;
razn_h_mem[8562] = 88;
razn_h_mem[8563] = 218;
razn_h_mem[8564] = 94;
razn_h_mem[8565] = 224;
razn_h_mem[8566] = 100;
razn_h_mem[8567] = 230;
razn_h_mem[8568] = 106;
razn_h_mem[8569] = 236;
razn_h_mem[8570] = 112;
razn_h_mem[8571] = 242;
razn_h_mem[8572] = 118;
razn_h_mem[8573] = 248;
razn_h_mem[8574] = 124;
razn_h_mem[8575] = 255;
razn_h_mem[8576] = 0;
razn_h_mem[8577] = 130;
razn_h_mem[8578] = 6;
razn_h_mem[8579] = 136;
razn_h_mem[8580] = 12;
razn_h_mem[8581] = 142;
razn_h_mem[8582] = 18;
razn_h_mem[8583] = 148;
razn_h_mem[8584] = 24;
razn_h_mem[8585] = 154;
razn_h_mem[8586] = 30;
razn_h_mem[8587] = 160;
razn_h_mem[8588] = 36;
razn_h_mem[8589] = 166;
razn_h_mem[8590] = 42;
razn_h_mem[8591] = 172;
razn_h_mem[8592] = 48;
razn_h_mem[8593] = 178;
razn_h_mem[8594] = 54;
razn_h_mem[8595] = 184;
razn_h_mem[8596] = 60;
razn_h_mem[8597] = 190;
razn_h_mem[8598] = 66;
razn_h_mem[8599] = 196;
razn_h_mem[8600] = 72;
razn_h_mem[8601] = 202;
razn_h_mem[8602] = 78;
razn_h_mem[8603] = 208;
razn_h_mem[8604] = 84;
razn_h_mem[8605] = 214;
razn_h_mem[8606] = 90;
razn_h_mem[8607] = 220;
razn_h_mem[8608] = 96;
razn_h_mem[8609] = 226;
razn_h_mem[8610] = 102;
razn_h_mem[8611] = 232;
razn_h_mem[8612] = 108;
razn_h_mem[8613] = 238;
razn_h_mem[8614] = 114;
razn_h_mem[8615] = 244;
razn_h_mem[8616] = 120;
razn_h_mem[8617] = 250;
razn_h_mem[8618] = 126;
razn_h_mem[8619] = 2;
razn_h_mem[8620] = 132;
razn_h_mem[8621] = 8;
razn_h_mem[8622] = 138;
razn_h_mem[8623] = 14;
razn_h_mem[8624] = 144;
razn_h_mem[8625] = 20;
razn_h_mem[8626] = 150;
razn_h_mem[8627] = 26;
razn_h_mem[8628] = 156;
razn_h_mem[8629] = 32;
razn_h_mem[8630] = 162;
razn_h_mem[8631] = 38;
razn_h_mem[8632] = 168;
razn_h_mem[8633] = 44;
razn_h_mem[8634] = 174;
razn_h_mem[8635] = 50;
razn_h_mem[8636] = 180;
razn_h_mem[8637] = 56;
razn_h_mem[8638] = 186;
razn_h_mem[8639] = 62;
razn_h_mem[8640] = 192;
razn_h_mem[8641] = 68;
razn_h_mem[8642] = 198;
razn_h_mem[8643] = 74;
razn_h_mem[8644] = 204;
razn_h_mem[8645] = 80;
razn_h_mem[8646] = 210;
razn_h_mem[8647] = 86;
razn_h_mem[8648] = 216;
razn_h_mem[8649] = 92;
razn_h_mem[8650] = 222;
razn_h_mem[8651] = 98;
razn_h_mem[8652] = 228;
razn_h_mem[8653] = 104;
razn_h_mem[8654] = 234;
razn_h_mem[8655] = 110;
razn_h_mem[8656] = 240;
razn_h_mem[8657] = 116;
razn_h_mem[8658] = 246;
razn_h_mem[8659] = 122;
razn_h_mem[8660] = 252;
razn_h_mem[8661] = 128;
razn_h_mem[8662] = 4;
razn_h_mem[8663] = 134;
razn_h_mem[8664] = 10;
razn_h_mem[8665] = 140;
razn_h_mem[8666] = 16;
razn_h_mem[8667] = 146;
razn_h_mem[8668] = 22;
razn_h_mem[8669] = 152;
razn_h_mem[8670] = 28;
razn_h_mem[8671] = 158;
razn_h_mem[8672] = 34;
razn_h_mem[8673] = 164;
razn_h_mem[8674] = 40;
razn_h_mem[8675] = 170;
razn_h_mem[8676] = 46;
razn_h_mem[8677] = 176;
razn_h_mem[8678] = 52;
razn_h_mem[8679] = 182;
razn_h_mem[8680] = 58;
razn_h_mem[8681] = 188;
razn_h_mem[8682] = 64;
razn_h_mem[8683] = 194;
razn_h_mem[8684] = 70;
razn_h_mem[8685] = 200;
razn_h_mem[8686] = 76;
razn_h_mem[8687] = 206;
razn_h_mem[8688] = 82;
razn_h_mem[8689] = 212;
razn_h_mem[8690] = 88;
razn_h_mem[8691] = 218;
razn_h_mem[8692] = 94;
razn_h_mem[8693] = 224;
razn_h_mem[8694] = 100;
razn_h_mem[8695] = 230;
razn_h_mem[8696] = 106;
razn_h_mem[8697] = 236;
razn_h_mem[8698] = 112;
razn_h_mem[8699] = 242;
razn_h_mem[8700] = 118;
razn_h_mem[8701] = 248;
razn_h_mem[8702] = 124;
razn_h_mem[8703] = 255;
razn_h_mem[8704] = 0;
razn_h_mem[8705] = 130;
razn_h_mem[8706] = 6;
razn_h_mem[8707] = 136;
razn_h_mem[8708] = 12;
razn_h_mem[8709] = 142;
razn_h_mem[8710] = 18;
razn_h_mem[8711] = 148;
razn_h_mem[8712] = 24;
razn_h_mem[8713] = 154;
razn_h_mem[8714] = 30;
razn_h_mem[8715] = 160;
razn_h_mem[8716] = 36;
razn_h_mem[8717] = 166;
razn_h_mem[8718] = 42;
razn_h_mem[8719] = 172;
razn_h_mem[8720] = 48;
razn_h_mem[8721] = 178;
razn_h_mem[8722] = 54;
razn_h_mem[8723] = 184;
razn_h_mem[8724] = 60;
razn_h_mem[8725] = 190;
razn_h_mem[8726] = 66;
razn_h_mem[8727] = 196;
razn_h_mem[8728] = 72;
razn_h_mem[8729] = 202;
razn_h_mem[8730] = 78;
razn_h_mem[8731] = 208;
razn_h_mem[8732] = 84;
razn_h_mem[8733] = 214;
razn_h_mem[8734] = 90;
razn_h_mem[8735] = 220;
razn_h_mem[8736] = 96;
razn_h_mem[8737] = 226;
razn_h_mem[8738] = 102;
razn_h_mem[8739] = 232;
razn_h_mem[8740] = 108;
razn_h_mem[8741] = 238;
razn_h_mem[8742] = 114;
razn_h_mem[8743] = 244;
razn_h_mem[8744] = 120;
razn_h_mem[8745] = 250;
razn_h_mem[8746] = 126;
razn_h_mem[8747] = 2;
razn_h_mem[8748] = 132;
razn_h_mem[8749] = 8;
razn_h_mem[8750] = 138;
razn_h_mem[8751] = 14;
razn_h_mem[8752] = 144;
razn_h_mem[8753] = 20;
razn_h_mem[8754] = 150;
razn_h_mem[8755] = 26;
razn_h_mem[8756] = 156;
razn_h_mem[8757] = 32;
razn_h_mem[8758] = 162;
razn_h_mem[8759] = 38;
razn_h_mem[8760] = 168;
razn_h_mem[8761] = 44;
razn_h_mem[8762] = 174;
razn_h_mem[8763] = 50;
razn_h_mem[8764] = 180;
razn_h_mem[8765] = 56;
razn_h_mem[8766] = 186;
razn_h_mem[8767] = 62;
razn_h_mem[8768] = 192;
razn_h_mem[8769] = 68;
razn_h_mem[8770] = 198;
razn_h_mem[8771] = 74;
razn_h_mem[8772] = 204;
razn_h_mem[8773] = 80;
razn_h_mem[8774] = 210;
razn_h_mem[8775] = 86;
razn_h_mem[8776] = 216;
razn_h_mem[8777] = 92;
razn_h_mem[8778] = 222;
razn_h_mem[8779] = 98;
razn_h_mem[8780] = 228;
razn_h_mem[8781] = 104;
razn_h_mem[8782] = 234;
razn_h_mem[8783] = 110;
razn_h_mem[8784] = 240;
razn_h_mem[8785] = 116;
razn_h_mem[8786] = 246;
razn_h_mem[8787] = 122;
razn_h_mem[8788] = 252;
razn_h_mem[8789] = 128;
razn_h_mem[8790] = 4;
razn_h_mem[8791] = 134;
razn_h_mem[8792] = 10;
razn_h_mem[8793] = 140;
razn_h_mem[8794] = 16;
razn_h_mem[8795] = 146;
razn_h_mem[8796] = 22;
razn_h_mem[8797] = 152;
razn_h_mem[8798] = 28;
razn_h_mem[8799] = 158;
razn_h_mem[8800] = 34;
razn_h_mem[8801] = 164;
razn_h_mem[8802] = 40;
razn_h_mem[8803] = 170;
razn_h_mem[8804] = 46;
razn_h_mem[8805] = 176;
razn_h_mem[8806] = 52;
razn_h_mem[8807] = 182;
razn_h_mem[8808] = 58;
razn_h_mem[8809] = 188;
razn_h_mem[8810] = 64;
razn_h_mem[8811] = 194;
razn_h_mem[8812] = 70;
razn_h_mem[8813] = 200;
razn_h_mem[8814] = 76;
razn_h_mem[8815] = 206;
razn_h_mem[8816] = 82;
razn_h_mem[8817] = 212;
razn_h_mem[8818] = 88;
razn_h_mem[8819] = 218;
razn_h_mem[8820] = 94;
razn_h_mem[8821] = 224;
razn_h_mem[8822] = 100;
razn_h_mem[8823] = 230;
razn_h_mem[8824] = 106;
razn_h_mem[8825] = 236;
razn_h_mem[8826] = 112;
razn_h_mem[8827] = 242;
razn_h_mem[8828] = 118;
razn_h_mem[8829] = 248;
razn_h_mem[8830] = 124;
razn_h_mem[8831] = 255;
razn_h_mem[8832] = 0;
razn_h_mem[8833] = 130;
razn_h_mem[8834] = 6;
razn_h_mem[8835] = 136;
razn_h_mem[8836] = 12;
razn_h_mem[8837] = 142;
razn_h_mem[8838] = 18;
razn_h_mem[8839] = 148;
razn_h_mem[8840] = 24;
razn_h_mem[8841] = 154;
razn_h_mem[8842] = 30;
razn_h_mem[8843] = 160;
razn_h_mem[8844] = 36;
razn_h_mem[8845] = 166;
razn_h_mem[8846] = 42;
razn_h_mem[8847] = 172;
razn_h_mem[8848] = 48;
razn_h_mem[8849] = 178;
razn_h_mem[8850] = 54;
razn_h_mem[8851] = 184;
razn_h_mem[8852] = 60;
razn_h_mem[8853] = 190;
razn_h_mem[8854] = 66;
razn_h_mem[8855] = 196;
razn_h_mem[8856] = 72;
razn_h_mem[8857] = 202;
razn_h_mem[8858] = 78;
razn_h_mem[8859] = 208;
razn_h_mem[8860] = 84;
razn_h_mem[8861] = 214;
razn_h_mem[8862] = 90;
razn_h_mem[8863] = 220;
razn_h_mem[8864] = 96;
razn_h_mem[8865] = 226;
razn_h_mem[8866] = 102;
razn_h_mem[8867] = 232;
razn_h_mem[8868] = 108;
razn_h_mem[8869] = 238;
razn_h_mem[8870] = 114;
razn_h_mem[8871] = 244;
razn_h_mem[8872] = 120;
razn_h_mem[8873] = 250;
razn_h_mem[8874] = 126;
razn_h_mem[8875] = 2;
razn_h_mem[8876] = 132;
razn_h_mem[8877] = 8;
razn_h_mem[8878] = 138;
razn_h_mem[8879] = 14;
razn_h_mem[8880] = 144;
razn_h_mem[8881] = 20;
razn_h_mem[8882] = 150;
razn_h_mem[8883] = 26;
razn_h_mem[8884] = 156;
razn_h_mem[8885] = 32;
razn_h_mem[8886] = 162;
razn_h_mem[8887] = 38;
razn_h_mem[8888] = 168;
razn_h_mem[8889] = 44;
razn_h_mem[8890] = 174;
razn_h_mem[8891] = 50;
razn_h_mem[8892] = 180;
razn_h_mem[8893] = 56;
razn_h_mem[8894] = 186;
razn_h_mem[8895] = 62;
razn_h_mem[8896] = 192;
razn_h_mem[8897] = 68;
razn_h_mem[8898] = 198;
razn_h_mem[8899] = 74;
razn_h_mem[8900] = 204;
razn_h_mem[8901] = 80;
razn_h_mem[8902] = 210;
razn_h_mem[8903] = 86;
razn_h_mem[8904] = 216;
razn_h_mem[8905] = 92;
razn_h_mem[8906] = 222;
razn_h_mem[8907] = 98;
razn_h_mem[8908] = 228;
razn_h_mem[8909] = 104;
razn_h_mem[8910] = 234;
razn_h_mem[8911] = 110;
razn_h_mem[8912] = 240;
razn_h_mem[8913] = 116;
razn_h_mem[8914] = 246;
razn_h_mem[8915] = 122;
razn_h_mem[8916] = 252;
razn_h_mem[8917] = 128;
razn_h_mem[8918] = 4;
razn_h_mem[8919] = 134;
razn_h_mem[8920] = 10;
razn_h_mem[8921] = 140;
razn_h_mem[8922] = 16;
razn_h_mem[8923] = 146;
razn_h_mem[8924] = 22;
razn_h_mem[8925] = 152;
razn_h_mem[8926] = 28;
razn_h_mem[8927] = 158;
razn_h_mem[8928] = 34;
razn_h_mem[8929] = 164;
razn_h_mem[8930] = 40;
razn_h_mem[8931] = 170;
razn_h_mem[8932] = 46;
razn_h_mem[8933] = 176;
razn_h_mem[8934] = 52;
razn_h_mem[8935] = 182;
razn_h_mem[8936] = 58;
razn_h_mem[8937] = 188;
razn_h_mem[8938] = 64;
razn_h_mem[8939] = 194;
razn_h_mem[8940] = 70;
razn_h_mem[8941] = 200;
razn_h_mem[8942] = 76;
razn_h_mem[8943] = 206;
razn_h_mem[8944] = 82;
razn_h_mem[8945] = 212;
razn_h_mem[8946] = 88;
razn_h_mem[8947] = 218;
razn_h_mem[8948] = 94;
razn_h_mem[8949] = 224;
razn_h_mem[8950] = 100;
razn_h_mem[8951] = 230;
razn_h_mem[8952] = 106;
razn_h_mem[8953] = 236;
razn_h_mem[8954] = 112;
razn_h_mem[8955] = 242;
razn_h_mem[8956] = 118;
razn_h_mem[8957] = 248;
razn_h_mem[8958] = 124;
razn_h_mem[8959] = 255;
razn_h_mem[8960] = 0;
razn_h_mem[8961] = 130;
razn_h_mem[8962] = 6;
razn_h_mem[8963] = 136;
razn_h_mem[8964] = 12;
razn_h_mem[8965] = 142;
razn_h_mem[8966] = 18;
razn_h_mem[8967] = 148;
razn_h_mem[8968] = 24;
razn_h_mem[8969] = 154;
razn_h_mem[8970] = 30;
razn_h_mem[8971] = 160;
razn_h_mem[8972] = 36;
razn_h_mem[8973] = 166;
razn_h_mem[8974] = 42;
razn_h_mem[8975] = 172;
razn_h_mem[8976] = 48;
razn_h_mem[8977] = 178;
razn_h_mem[8978] = 54;
razn_h_mem[8979] = 184;
razn_h_mem[8980] = 60;
razn_h_mem[8981] = 190;
razn_h_mem[8982] = 66;
razn_h_mem[8983] = 196;
razn_h_mem[8984] = 72;
razn_h_mem[8985] = 202;
razn_h_mem[8986] = 78;
razn_h_mem[8987] = 208;
razn_h_mem[8988] = 84;
razn_h_mem[8989] = 214;
razn_h_mem[8990] = 90;
razn_h_mem[8991] = 220;
razn_h_mem[8992] = 96;
razn_h_mem[8993] = 226;
razn_h_mem[8994] = 102;
razn_h_mem[8995] = 232;
razn_h_mem[8996] = 108;
razn_h_mem[8997] = 238;
razn_h_mem[8998] = 114;
razn_h_mem[8999] = 244;
razn_h_mem[9000] = 120;
razn_h_mem[9001] = 250;
razn_h_mem[9002] = 126;
razn_h_mem[9003] = 2;
razn_h_mem[9004] = 132;
razn_h_mem[9005] = 8;
razn_h_mem[9006] = 138;
razn_h_mem[9007] = 14;
razn_h_mem[9008] = 144;
razn_h_mem[9009] = 20;
razn_h_mem[9010] = 150;
razn_h_mem[9011] = 26;
razn_h_mem[9012] = 156;
razn_h_mem[9013] = 32;
razn_h_mem[9014] = 162;
razn_h_mem[9015] = 38;
razn_h_mem[9016] = 168;
razn_h_mem[9017] = 44;
razn_h_mem[9018] = 174;
razn_h_mem[9019] = 50;
razn_h_mem[9020] = 180;
razn_h_mem[9021] = 56;
razn_h_mem[9022] = 186;
razn_h_mem[9023] = 62;
razn_h_mem[9024] = 192;
razn_h_mem[9025] = 68;
razn_h_mem[9026] = 198;
razn_h_mem[9027] = 74;
razn_h_mem[9028] = 204;
razn_h_mem[9029] = 80;
razn_h_mem[9030] = 210;
razn_h_mem[9031] = 86;
razn_h_mem[9032] = 216;
razn_h_mem[9033] = 92;
razn_h_mem[9034] = 222;
razn_h_mem[9035] = 98;
razn_h_mem[9036] = 228;
razn_h_mem[9037] = 104;
razn_h_mem[9038] = 234;
razn_h_mem[9039] = 110;
razn_h_mem[9040] = 240;
razn_h_mem[9041] = 116;
razn_h_mem[9042] = 246;
razn_h_mem[9043] = 122;
razn_h_mem[9044] = 252;
razn_h_mem[9045] = 128;
razn_h_mem[9046] = 4;
razn_h_mem[9047] = 134;
razn_h_mem[9048] = 10;
razn_h_mem[9049] = 140;
razn_h_mem[9050] = 16;
razn_h_mem[9051] = 146;
razn_h_mem[9052] = 22;
razn_h_mem[9053] = 152;
razn_h_mem[9054] = 28;
razn_h_mem[9055] = 158;
razn_h_mem[9056] = 34;
razn_h_mem[9057] = 164;
razn_h_mem[9058] = 40;
razn_h_mem[9059] = 170;
razn_h_mem[9060] = 46;
razn_h_mem[9061] = 176;
razn_h_mem[9062] = 52;
razn_h_mem[9063] = 182;
razn_h_mem[9064] = 58;
razn_h_mem[9065] = 188;
razn_h_mem[9066] = 64;
razn_h_mem[9067] = 194;
razn_h_mem[9068] = 70;
razn_h_mem[9069] = 200;
razn_h_mem[9070] = 76;
razn_h_mem[9071] = 206;
razn_h_mem[9072] = 82;
razn_h_mem[9073] = 212;
razn_h_mem[9074] = 88;
razn_h_mem[9075] = 218;
razn_h_mem[9076] = 94;
razn_h_mem[9077] = 224;
razn_h_mem[9078] = 100;
razn_h_mem[9079] = 230;
razn_h_mem[9080] = 106;
razn_h_mem[9081] = 236;
razn_h_mem[9082] = 112;
razn_h_mem[9083] = 242;
razn_h_mem[9084] = 118;
razn_h_mem[9085] = 248;
razn_h_mem[9086] = 124;
razn_h_mem[9087] = 255;
razn_h_mem[9088] = 0;
razn_h_mem[9089] = 130;
razn_h_mem[9090] = 6;
razn_h_mem[9091] = 136;
razn_h_mem[9092] = 12;
razn_h_mem[9093] = 142;
razn_h_mem[9094] = 18;
razn_h_mem[9095] = 148;
razn_h_mem[9096] = 24;
razn_h_mem[9097] = 154;
razn_h_mem[9098] = 30;
razn_h_mem[9099] = 160;
razn_h_mem[9100] = 36;
razn_h_mem[9101] = 166;
razn_h_mem[9102] = 42;
razn_h_mem[9103] = 172;
razn_h_mem[9104] = 48;
razn_h_mem[9105] = 178;
razn_h_mem[9106] = 54;
razn_h_mem[9107] = 184;
razn_h_mem[9108] = 60;
razn_h_mem[9109] = 190;
razn_h_mem[9110] = 66;
razn_h_mem[9111] = 196;
razn_h_mem[9112] = 72;
razn_h_mem[9113] = 202;
razn_h_mem[9114] = 78;
razn_h_mem[9115] = 208;
razn_h_mem[9116] = 84;
razn_h_mem[9117] = 214;
razn_h_mem[9118] = 90;
razn_h_mem[9119] = 220;
razn_h_mem[9120] = 96;
razn_h_mem[9121] = 226;
razn_h_mem[9122] = 102;
razn_h_mem[9123] = 232;
razn_h_mem[9124] = 108;
razn_h_mem[9125] = 238;
razn_h_mem[9126] = 114;
razn_h_mem[9127] = 244;
razn_h_mem[9128] = 120;
razn_h_mem[9129] = 250;
razn_h_mem[9130] = 126;
razn_h_mem[9131] = 2;
razn_h_mem[9132] = 132;
razn_h_mem[9133] = 8;
razn_h_mem[9134] = 138;
razn_h_mem[9135] = 14;
razn_h_mem[9136] = 144;
razn_h_mem[9137] = 20;
razn_h_mem[9138] = 150;
razn_h_mem[9139] = 26;
razn_h_mem[9140] = 156;
razn_h_mem[9141] = 32;
razn_h_mem[9142] = 162;
razn_h_mem[9143] = 38;
razn_h_mem[9144] = 168;
razn_h_mem[9145] = 44;
razn_h_mem[9146] = 174;
razn_h_mem[9147] = 50;
razn_h_mem[9148] = 180;
razn_h_mem[9149] = 56;
razn_h_mem[9150] = 186;
razn_h_mem[9151] = 62;
razn_h_mem[9152] = 192;
razn_h_mem[9153] = 68;
razn_h_mem[9154] = 198;
razn_h_mem[9155] = 74;
razn_h_mem[9156] = 204;
razn_h_mem[9157] = 80;
razn_h_mem[9158] = 210;
razn_h_mem[9159] = 86;
razn_h_mem[9160] = 216;
razn_h_mem[9161] = 92;
razn_h_mem[9162] = 222;
razn_h_mem[9163] = 98;
razn_h_mem[9164] = 228;
razn_h_mem[9165] = 104;
razn_h_mem[9166] = 234;
razn_h_mem[9167] = 110;
razn_h_mem[9168] = 240;
razn_h_mem[9169] = 116;
razn_h_mem[9170] = 246;
razn_h_mem[9171] = 122;
razn_h_mem[9172] = 252;
razn_h_mem[9173] = 128;
razn_h_mem[9174] = 4;
razn_h_mem[9175] = 134;
razn_h_mem[9176] = 10;
razn_h_mem[9177] = 140;
razn_h_mem[9178] = 16;
razn_h_mem[9179] = 146;
razn_h_mem[9180] = 22;
razn_h_mem[9181] = 152;
razn_h_mem[9182] = 28;
razn_h_mem[9183] = 158;
razn_h_mem[9184] = 34;
razn_h_mem[9185] = 164;
razn_h_mem[9186] = 40;
razn_h_mem[9187] = 170;
razn_h_mem[9188] = 46;
razn_h_mem[9189] = 176;
razn_h_mem[9190] = 52;
razn_h_mem[9191] = 182;
razn_h_mem[9192] = 58;
razn_h_mem[9193] = 188;
razn_h_mem[9194] = 64;
razn_h_mem[9195] = 194;
razn_h_mem[9196] = 70;
razn_h_mem[9197] = 200;
razn_h_mem[9198] = 76;
razn_h_mem[9199] = 206;
razn_h_mem[9200] = 82;
razn_h_mem[9201] = 212;
razn_h_mem[9202] = 88;
razn_h_mem[9203] = 218;
razn_h_mem[9204] = 94;
razn_h_mem[9205] = 224;
razn_h_mem[9206] = 100;
razn_h_mem[9207] = 230;
razn_h_mem[9208] = 106;
razn_h_mem[9209] = 236;
razn_h_mem[9210] = 112;
razn_h_mem[9211] = 242;
razn_h_mem[9212] = 118;
razn_h_mem[9213] = 248;
razn_h_mem[9214] = 124;
razn_h_mem[9215] = 255;
razn_h_mem[9216] = 0;
razn_h_mem[9217] = 130;
razn_h_mem[9218] = 6;
razn_h_mem[9219] = 136;
razn_h_mem[9220] = 12;
razn_h_mem[9221] = 142;
razn_h_mem[9222] = 18;
razn_h_mem[9223] = 148;
razn_h_mem[9224] = 24;
razn_h_mem[9225] = 154;
razn_h_mem[9226] = 30;
razn_h_mem[9227] = 160;
razn_h_mem[9228] = 36;
razn_h_mem[9229] = 166;
razn_h_mem[9230] = 42;
razn_h_mem[9231] = 172;
razn_h_mem[9232] = 48;
razn_h_mem[9233] = 178;
razn_h_mem[9234] = 54;
razn_h_mem[9235] = 184;
razn_h_mem[9236] = 60;
razn_h_mem[9237] = 190;
razn_h_mem[9238] = 66;
razn_h_mem[9239] = 196;
razn_h_mem[9240] = 72;
razn_h_mem[9241] = 202;
razn_h_mem[9242] = 78;
razn_h_mem[9243] = 208;
razn_h_mem[9244] = 84;
razn_h_mem[9245] = 214;
razn_h_mem[9246] = 90;
razn_h_mem[9247] = 220;
razn_h_mem[9248] = 96;
razn_h_mem[9249] = 226;
razn_h_mem[9250] = 102;
razn_h_mem[9251] = 232;
razn_h_mem[9252] = 108;
razn_h_mem[9253] = 238;
razn_h_mem[9254] = 114;
razn_h_mem[9255] = 244;
razn_h_mem[9256] = 120;
razn_h_mem[9257] = 250;
razn_h_mem[9258] = 126;
razn_h_mem[9259] = 2;
razn_h_mem[9260] = 132;
razn_h_mem[9261] = 8;
razn_h_mem[9262] = 138;
razn_h_mem[9263] = 14;
razn_h_mem[9264] = 144;
razn_h_mem[9265] = 20;
razn_h_mem[9266] = 150;
razn_h_mem[9267] = 26;
razn_h_mem[9268] = 156;
razn_h_mem[9269] = 32;
razn_h_mem[9270] = 162;
razn_h_mem[9271] = 38;
razn_h_mem[9272] = 168;
razn_h_mem[9273] = 44;
razn_h_mem[9274] = 174;
razn_h_mem[9275] = 50;
razn_h_mem[9276] = 180;
razn_h_mem[9277] = 56;
razn_h_mem[9278] = 186;
razn_h_mem[9279] = 62;
razn_h_mem[9280] = 192;
razn_h_mem[9281] = 68;
razn_h_mem[9282] = 198;
razn_h_mem[9283] = 74;
razn_h_mem[9284] = 204;
razn_h_mem[9285] = 80;
razn_h_mem[9286] = 210;
razn_h_mem[9287] = 86;
razn_h_mem[9288] = 216;
razn_h_mem[9289] = 92;
razn_h_mem[9290] = 222;
razn_h_mem[9291] = 98;
razn_h_mem[9292] = 228;
razn_h_mem[9293] = 104;
razn_h_mem[9294] = 234;
razn_h_mem[9295] = 110;
razn_h_mem[9296] = 240;
razn_h_mem[9297] = 116;
razn_h_mem[9298] = 246;
razn_h_mem[9299] = 122;
razn_h_mem[9300] = 252;
razn_h_mem[9301] = 128;
razn_h_mem[9302] = 4;
razn_h_mem[9303] = 134;
razn_h_mem[9304] = 10;
razn_h_mem[9305] = 140;
razn_h_mem[9306] = 16;
razn_h_mem[9307] = 146;
razn_h_mem[9308] = 22;
razn_h_mem[9309] = 152;
razn_h_mem[9310] = 28;
razn_h_mem[9311] = 158;
razn_h_mem[9312] = 34;
razn_h_mem[9313] = 164;
razn_h_mem[9314] = 40;
razn_h_mem[9315] = 170;
razn_h_mem[9316] = 46;
razn_h_mem[9317] = 176;
razn_h_mem[9318] = 52;
razn_h_mem[9319] = 182;
razn_h_mem[9320] = 58;
razn_h_mem[9321] = 188;
razn_h_mem[9322] = 64;
razn_h_mem[9323] = 194;
razn_h_mem[9324] = 70;
razn_h_mem[9325] = 200;
razn_h_mem[9326] = 76;
razn_h_mem[9327] = 206;
razn_h_mem[9328] = 82;
razn_h_mem[9329] = 212;
razn_h_mem[9330] = 88;
razn_h_mem[9331] = 218;
razn_h_mem[9332] = 94;
razn_h_mem[9333] = 224;
razn_h_mem[9334] = 100;
razn_h_mem[9335] = 230;
razn_h_mem[9336] = 106;
razn_h_mem[9337] = 236;
razn_h_mem[9338] = 112;
razn_h_mem[9339] = 242;
razn_h_mem[9340] = 118;
razn_h_mem[9341] = 248;
razn_h_mem[9342] = 124;
razn_h_mem[9343] = 255;
razn_h_mem[9344] = 0;
razn_h_mem[9345] = 130;
razn_h_mem[9346] = 6;
razn_h_mem[9347] = 136;
razn_h_mem[9348] = 12;
razn_h_mem[9349] = 142;
razn_h_mem[9350] = 18;
razn_h_mem[9351] = 148;
razn_h_mem[9352] = 24;
razn_h_mem[9353] = 154;
razn_h_mem[9354] = 30;
razn_h_mem[9355] = 160;
razn_h_mem[9356] = 36;
razn_h_mem[9357] = 166;
razn_h_mem[9358] = 42;
razn_h_mem[9359] = 172;
razn_h_mem[9360] = 48;
razn_h_mem[9361] = 178;
razn_h_mem[9362] = 54;
razn_h_mem[9363] = 184;
razn_h_mem[9364] = 60;
razn_h_mem[9365] = 190;
razn_h_mem[9366] = 66;
razn_h_mem[9367] = 196;
razn_h_mem[9368] = 72;
razn_h_mem[9369] = 202;
razn_h_mem[9370] = 78;
razn_h_mem[9371] = 208;
razn_h_mem[9372] = 84;
razn_h_mem[9373] = 214;
razn_h_mem[9374] = 90;
razn_h_mem[9375] = 220;
razn_h_mem[9376] = 96;
razn_h_mem[9377] = 226;
razn_h_mem[9378] = 102;
razn_h_mem[9379] = 232;
razn_h_mem[9380] = 108;
razn_h_mem[9381] = 238;
razn_h_mem[9382] = 114;
razn_h_mem[9383] = 244;
razn_h_mem[9384] = 120;
razn_h_mem[9385] = 250;
razn_h_mem[9386] = 126;
razn_h_mem[9387] = 2;
razn_h_mem[9388] = 132;
razn_h_mem[9389] = 8;
razn_h_mem[9390] = 138;
razn_h_mem[9391] = 14;
razn_h_mem[9392] = 144;
razn_h_mem[9393] = 20;
razn_h_mem[9394] = 150;
razn_h_mem[9395] = 26;
razn_h_mem[9396] = 156;
razn_h_mem[9397] = 32;
razn_h_mem[9398] = 162;
razn_h_mem[9399] = 38;
razn_h_mem[9400] = 168;
razn_h_mem[9401] = 44;
razn_h_mem[9402] = 174;
razn_h_mem[9403] = 50;
razn_h_mem[9404] = 180;
razn_h_mem[9405] = 56;
razn_h_mem[9406] = 186;
razn_h_mem[9407] = 62;
razn_h_mem[9408] = 192;
razn_h_mem[9409] = 68;
razn_h_mem[9410] = 198;
razn_h_mem[9411] = 74;
razn_h_mem[9412] = 204;
razn_h_mem[9413] = 80;
razn_h_mem[9414] = 210;
razn_h_mem[9415] = 86;
razn_h_mem[9416] = 216;
razn_h_mem[9417] = 92;
razn_h_mem[9418] = 222;
razn_h_mem[9419] = 98;
razn_h_mem[9420] = 228;
razn_h_mem[9421] = 104;
razn_h_mem[9422] = 234;
razn_h_mem[9423] = 110;
razn_h_mem[9424] = 240;
razn_h_mem[9425] = 116;
razn_h_mem[9426] = 246;
razn_h_mem[9427] = 122;
razn_h_mem[9428] = 252;
razn_h_mem[9429] = 128;
razn_h_mem[9430] = 4;
razn_h_mem[9431] = 134;
razn_h_mem[9432] = 10;
razn_h_mem[9433] = 140;
razn_h_mem[9434] = 16;
razn_h_mem[9435] = 146;
razn_h_mem[9436] = 22;
razn_h_mem[9437] = 152;
razn_h_mem[9438] = 28;
razn_h_mem[9439] = 158;
razn_h_mem[9440] = 34;
razn_h_mem[9441] = 164;
razn_h_mem[9442] = 40;
razn_h_mem[9443] = 170;
razn_h_mem[9444] = 46;
razn_h_mem[9445] = 176;
razn_h_mem[9446] = 52;
razn_h_mem[9447] = 182;
razn_h_mem[9448] = 58;
razn_h_mem[9449] = 188;
razn_h_mem[9450] = 64;
razn_h_mem[9451] = 194;
razn_h_mem[9452] = 70;
razn_h_mem[9453] = 200;
razn_h_mem[9454] = 76;
razn_h_mem[9455] = 206;
razn_h_mem[9456] = 82;
razn_h_mem[9457] = 212;
razn_h_mem[9458] = 88;
razn_h_mem[9459] = 218;
razn_h_mem[9460] = 94;
razn_h_mem[9461] = 224;
razn_h_mem[9462] = 100;
razn_h_mem[9463] = 230;
razn_h_mem[9464] = 106;
razn_h_mem[9465] = 236;
razn_h_mem[9466] = 112;
razn_h_mem[9467] = 242;
razn_h_mem[9468] = 118;
razn_h_mem[9469] = 248;
razn_h_mem[9470] = 124;
razn_h_mem[9471] = 255;
razn_h_mem[9472] = 0;
razn_h_mem[9473] = 130;
razn_h_mem[9474] = 6;
razn_h_mem[9475] = 136;
razn_h_mem[9476] = 12;
razn_h_mem[9477] = 142;
razn_h_mem[9478] = 18;
razn_h_mem[9479] = 148;
razn_h_mem[9480] = 24;
razn_h_mem[9481] = 154;
razn_h_mem[9482] = 30;
razn_h_mem[9483] = 160;
razn_h_mem[9484] = 36;
razn_h_mem[9485] = 166;
razn_h_mem[9486] = 42;
razn_h_mem[9487] = 172;
razn_h_mem[9488] = 48;
razn_h_mem[9489] = 178;
razn_h_mem[9490] = 54;
razn_h_mem[9491] = 184;
razn_h_mem[9492] = 60;
razn_h_mem[9493] = 190;
razn_h_mem[9494] = 66;
razn_h_mem[9495] = 196;
razn_h_mem[9496] = 72;
razn_h_mem[9497] = 202;
razn_h_mem[9498] = 78;
razn_h_mem[9499] = 208;
razn_h_mem[9500] = 84;
razn_h_mem[9501] = 214;
razn_h_mem[9502] = 90;
razn_h_mem[9503] = 220;
razn_h_mem[9504] = 96;
razn_h_mem[9505] = 226;
razn_h_mem[9506] = 102;
razn_h_mem[9507] = 232;
razn_h_mem[9508] = 108;
razn_h_mem[9509] = 238;
razn_h_mem[9510] = 114;
razn_h_mem[9511] = 244;
razn_h_mem[9512] = 120;
razn_h_mem[9513] = 250;
razn_h_mem[9514] = 126;
razn_h_mem[9515] = 2;
razn_h_mem[9516] = 132;
razn_h_mem[9517] = 8;
razn_h_mem[9518] = 138;
razn_h_mem[9519] = 14;
razn_h_mem[9520] = 144;
razn_h_mem[9521] = 20;
razn_h_mem[9522] = 150;
razn_h_mem[9523] = 26;
razn_h_mem[9524] = 156;
razn_h_mem[9525] = 32;
razn_h_mem[9526] = 162;
razn_h_mem[9527] = 38;
razn_h_mem[9528] = 168;
razn_h_mem[9529] = 44;
razn_h_mem[9530] = 174;
razn_h_mem[9531] = 50;
razn_h_mem[9532] = 180;
razn_h_mem[9533] = 56;
razn_h_mem[9534] = 186;
razn_h_mem[9535] = 62;
razn_h_mem[9536] = 192;
razn_h_mem[9537] = 68;
razn_h_mem[9538] = 198;
razn_h_mem[9539] = 74;
razn_h_mem[9540] = 204;
razn_h_mem[9541] = 80;
razn_h_mem[9542] = 210;
razn_h_mem[9543] = 86;
razn_h_mem[9544] = 216;
razn_h_mem[9545] = 92;
razn_h_mem[9546] = 222;
razn_h_mem[9547] = 98;
razn_h_mem[9548] = 228;
razn_h_mem[9549] = 104;
razn_h_mem[9550] = 234;
razn_h_mem[9551] = 110;
razn_h_mem[9552] = 240;
razn_h_mem[9553] = 116;
razn_h_mem[9554] = 246;
razn_h_mem[9555] = 122;
razn_h_mem[9556] = 252;
razn_h_mem[9557] = 128;
razn_h_mem[9558] = 4;
razn_h_mem[9559] = 134;
razn_h_mem[9560] = 10;
razn_h_mem[9561] = 140;
razn_h_mem[9562] = 16;
razn_h_mem[9563] = 146;
razn_h_mem[9564] = 22;
razn_h_mem[9565] = 152;
razn_h_mem[9566] = 28;
razn_h_mem[9567] = 158;
razn_h_mem[9568] = 34;
razn_h_mem[9569] = 164;
razn_h_mem[9570] = 40;
razn_h_mem[9571] = 170;
razn_h_mem[9572] = 46;
razn_h_mem[9573] = 176;
razn_h_mem[9574] = 52;
razn_h_mem[9575] = 182;
razn_h_mem[9576] = 58;
razn_h_mem[9577] = 188;
razn_h_mem[9578] = 64;
razn_h_mem[9579] = 194;
razn_h_mem[9580] = 70;
razn_h_mem[9581] = 200;
razn_h_mem[9582] = 76;
razn_h_mem[9583] = 206;
razn_h_mem[9584] = 82;
razn_h_mem[9585] = 212;
razn_h_mem[9586] = 88;
razn_h_mem[9587] = 218;
razn_h_mem[9588] = 94;
razn_h_mem[9589] = 224;
razn_h_mem[9590] = 100;
razn_h_mem[9591] = 230;
razn_h_mem[9592] = 106;
razn_h_mem[9593] = 236;
razn_h_mem[9594] = 112;
razn_h_mem[9595] = 242;
razn_h_mem[9596] = 118;
razn_h_mem[9597] = 248;
razn_h_mem[9598] = 124;
razn_h_mem[9599] = 255;
razn_h_mem[9600] = 0;
razn_h_mem[9601] = 130;
razn_h_mem[9602] = 6;
razn_h_mem[9603] = 136;
razn_h_mem[9604] = 12;
razn_h_mem[9605] = 142;
razn_h_mem[9606] = 18;
razn_h_mem[9607] = 148;
razn_h_mem[9608] = 24;
razn_h_mem[9609] = 154;
razn_h_mem[9610] = 30;
razn_h_mem[9611] = 160;
razn_h_mem[9612] = 36;
razn_h_mem[9613] = 166;
razn_h_mem[9614] = 42;
razn_h_mem[9615] = 172;
razn_h_mem[9616] = 48;
razn_h_mem[9617] = 178;
razn_h_mem[9618] = 54;
razn_h_mem[9619] = 184;
razn_h_mem[9620] = 60;
razn_h_mem[9621] = 190;
razn_h_mem[9622] = 66;
razn_h_mem[9623] = 196;
razn_h_mem[9624] = 72;
razn_h_mem[9625] = 202;
razn_h_mem[9626] = 78;
razn_h_mem[9627] = 208;
razn_h_mem[9628] = 84;
razn_h_mem[9629] = 214;
razn_h_mem[9630] = 90;
razn_h_mem[9631] = 220;
razn_h_mem[9632] = 96;
razn_h_mem[9633] = 226;
razn_h_mem[9634] = 102;
razn_h_mem[9635] = 232;
razn_h_mem[9636] = 108;
razn_h_mem[9637] = 238;
razn_h_mem[9638] = 114;
razn_h_mem[9639] = 244;
razn_h_mem[9640] = 120;
razn_h_mem[9641] = 250;
razn_h_mem[9642] = 126;
razn_h_mem[9643] = 2;
razn_h_mem[9644] = 132;
razn_h_mem[9645] = 8;
razn_h_mem[9646] = 138;
razn_h_mem[9647] = 14;
razn_h_mem[9648] = 144;
razn_h_mem[9649] = 20;
razn_h_mem[9650] = 150;
razn_h_mem[9651] = 26;
razn_h_mem[9652] = 156;
razn_h_mem[9653] = 32;
razn_h_mem[9654] = 162;
razn_h_mem[9655] = 38;
razn_h_mem[9656] = 168;
razn_h_mem[9657] = 44;
razn_h_mem[9658] = 174;
razn_h_mem[9659] = 50;
razn_h_mem[9660] = 180;
razn_h_mem[9661] = 56;
razn_h_mem[9662] = 186;
razn_h_mem[9663] = 62;
razn_h_mem[9664] = 192;
razn_h_mem[9665] = 68;
razn_h_mem[9666] = 198;
razn_h_mem[9667] = 74;
razn_h_mem[9668] = 204;
razn_h_mem[9669] = 80;
razn_h_mem[9670] = 210;
razn_h_mem[9671] = 86;
razn_h_mem[9672] = 216;
razn_h_mem[9673] = 92;
razn_h_mem[9674] = 222;
razn_h_mem[9675] = 98;
razn_h_mem[9676] = 228;
razn_h_mem[9677] = 104;
razn_h_mem[9678] = 234;
razn_h_mem[9679] = 110;
razn_h_mem[9680] = 240;
razn_h_mem[9681] = 116;
razn_h_mem[9682] = 246;
razn_h_mem[9683] = 122;
razn_h_mem[9684] = 252;
razn_h_mem[9685] = 128;
razn_h_mem[9686] = 4;
razn_h_mem[9687] = 134;
razn_h_mem[9688] = 10;
razn_h_mem[9689] = 140;
razn_h_mem[9690] = 16;
razn_h_mem[9691] = 146;
razn_h_mem[9692] = 22;
razn_h_mem[9693] = 152;
razn_h_mem[9694] = 28;
razn_h_mem[9695] = 158;
razn_h_mem[9696] = 34;
razn_h_mem[9697] = 164;
razn_h_mem[9698] = 40;
razn_h_mem[9699] = 170;
razn_h_mem[9700] = 46;
razn_h_mem[9701] = 176;
razn_h_mem[9702] = 52;
razn_h_mem[9703] = 182;
razn_h_mem[9704] = 58;
razn_h_mem[9705] = 188;
razn_h_mem[9706] = 64;
razn_h_mem[9707] = 194;
razn_h_mem[9708] = 70;
razn_h_mem[9709] = 200;
razn_h_mem[9710] = 76;
razn_h_mem[9711] = 206;
razn_h_mem[9712] = 82;
razn_h_mem[9713] = 212;
razn_h_mem[9714] = 88;
razn_h_mem[9715] = 218;
razn_h_mem[9716] = 94;
razn_h_mem[9717] = 224;
razn_h_mem[9718] = 100;
razn_h_mem[9719] = 230;
razn_h_mem[9720] = 106;
razn_h_mem[9721] = 236;
razn_h_mem[9722] = 112;
razn_h_mem[9723] = 242;
razn_h_mem[9724] = 118;
razn_h_mem[9725] = 248;
razn_h_mem[9726] = 124;
razn_h_mem[9727] = 255;
razn_h_mem[9728] = 0;
razn_h_mem[9729] = 130;
razn_h_mem[9730] = 6;
razn_h_mem[9731] = 136;
razn_h_mem[9732] = 12;
razn_h_mem[9733] = 142;
razn_h_mem[9734] = 18;
razn_h_mem[9735] = 148;
razn_h_mem[9736] = 24;
razn_h_mem[9737] = 154;
razn_h_mem[9738] = 30;
razn_h_mem[9739] = 160;
razn_h_mem[9740] = 36;
razn_h_mem[9741] = 166;
razn_h_mem[9742] = 42;
razn_h_mem[9743] = 172;
razn_h_mem[9744] = 48;
razn_h_mem[9745] = 178;
razn_h_mem[9746] = 54;
razn_h_mem[9747] = 184;
razn_h_mem[9748] = 60;
razn_h_mem[9749] = 190;
razn_h_mem[9750] = 66;
razn_h_mem[9751] = 196;
razn_h_mem[9752] = 72;
razn_h_mem[9753] = 202;
razn_h_mem[9754] = 78;
razn_h_mem[9755] = 208;
razn_h_mem[9756] = 84;
razn_h_mem[9757] = 214;
razn_h_mem[9758] = 90;
razn_h_mem[9759] = 220;
razn_h_mem[9760] = 96;
razn_h_mem[9761] = 226;
razn_h_mem[9762] = 102;
razn_h_mem[9763] = 232;
razn_h_mem[9764] = 108;
razn_h_mem[9765] = 238;
razn_h_mem[9766] = 114;
razn_h_mem[9767] = 244;
razn_h_mem[9768] = 120;
razn_h_mem[9769] = 250;
razn_h_mem[9770] = 126;
razn_h_mem[9771] = 2;
razn_h_mem[9772] = 132;
razn_h_mem[9773] = 8;
razn_h_mem[9774] = 138;
razn_h_mem[9775] = 14;
razn_h_mem[9776] = 144;
razn_h_mem[9777] = 20;
razn_h_mem[9778] = 150;
razn_h_mem[9779] = 26;
razn_h_mem[9780] = 156;
razn_h_mem[9781] = 32;
razn_h_mem[9782] = 162;
razn_h_mem[9783] = 38;
razn_h_mem[9784] = 168;
razn_h_mem[9785] = 44;
razn_h_mem[9786] = 174;
razn_h_mem[9787] = 50;
razn_h_mem[9788] = 180;
razn_h_mem[9789] = 56;
razn_h_mem[9790] = 186;
razn_h_mem[9791] = 62;
razn_h_mem[9792] = 192;
razn_h_mem[9793] = 68;
razn_h_mem[9794] = 198;
razn_h_mem[9795] = 74;
razn_h_mem[9796] = 204;
razn_h_mem[9797] = 80;
razn_h_mem[9798] = 210;
razn_h_mem[9799] = 86;
razn_h_mem[9800] = 216;
razn_h_mem[9801] = 92;
razn_h_mem[9802] = 222;
razn_h_mem[9803] = 98;
razn_h_mem[9804] = 228;
razn_h_mem[9805] = 104;
razn_h_mem[9806] = 234;
razn_h_mem[9807] = 110;
razn_h_mem[9808] = 240;
razn_h_mem[9809] = 116;
razn_h_mem[9810] = 246;
razn_h_mem[9811] = 122;
razn_h_mem[9812] = 252;
razn_h_mem[9813] = 128;
razn_h_mem[9814] = 4;
razn_h_mem[9815] = 134;
razn_h_mem[9816] = 10;
razn_h_mem[9817] = 140;
razn_h_mem[9818] = 16;
razn_h_mem[9819] = 146;
razn_h_mem[9820] = 22;
razn_h_mem[9821] = 152;
razn_h_mem[9822] = 28;
razn_h_mem[9823] = 158;
razn_h_mem[9824] = 34;
razn_h_mem[9825] = 164;
razn_h_mem[9826] = 40;
razn_h_mem[9827] = 170;
razn_h_mem[9828] = 46;
razn_h_mem[9829] = 176;
razn_h_mem[9830] = 52;
razn_h_mem[9831] = 182;
razn_h_mem[9832] = 58;
razn_h_mem[9833] = 188;
razn_h_mem[9834] = 64;
razn_h_mem[9835] = 194;
razn_h_mem[9836] = 70;
razn_h_mem[9837] = 200;
razn_h_mem[9838] = 76;
razn_h_mem[9839] = 206;
razn_h_mem[9840] = 82;
razn_h_mem[9841] = 212;
razn_h_mem[9842] = 88;
razn_h_mem[9843] = 218;
razn_h_mem[9844] = 94;
razn_h_mem[9845] = 224;
razn_h_mem[9846] = 100;
razn_h_mem[9847] = 230;
razn_h_mem[9848] = 106;
razn_h_mem[9849] = 236;
razn_h_mem[9850] = 112;
razn_h_mem[9851] = 242;
razn_h_mem[9852] = 118;
razn_h_mem[9853] = 248;
razn_h_mem[9854] = 124;
razn_h_mem[9855] = 255;
razn_h_mem[9856] = 0;
razn_h_mem[9857] = 130;
razn_h_mem[9858] = 6;
razn_h_mem[9859] = 136;
razn_h_mem[9860] = 12;
razn_h_mem[9861] = 142;
razn_h_mem[9862] = 18;
razn_h_mem[9863] = 148;
razn_h_mem[9864] = 24;
razn_h_mem[9865] = 154;
razn_h_mem[9866] = 30;
razn_h_mem[9867] = 160;
razn_h_mem[9868] = 36;
razn_h_mem[9869] = 166;
razn_h_mem[9870] = 42;
razn_h_mem[9871] = 172;
razn_h_mem[9872] = 48;
razn_h_mem[9873] = 178;
razn_h_mem[9874] = 54;
razn_h_mem[9875] = 184;
razn_h_mem[9876] = 60;
razn_h_mem[9877] = 190;
razn_h_mem[9878] = 66;
razn_h_mem[9879] = 196;
razn_h_mem[9880] = 72;
razn_h_mem[9881] = 202;
razn_h_mem[9882] = 78;
razn_h_mem[9883] = 208;
razn_h_mem[9884] = 84;
razn_h_mem[9885] = 214;
razn_h_mem[9886] = 90;
razn_h_mem[9887] = 220;
razn_h_mem[9888] = 96;
razn_h_mem[9889] = 226;
razn_h_mem[9890] = 102;
razn_h_mem[9891] = 232;
razn_h_mem[9892] = 108;
razn_h_mem[9893] = 238;
razn_h_mem[9894] = 114;
razn_h_mem[9895] = 244;
razn_h_mem[9896] = 120;
razn_h_mem[9897] = 250;
razn_h_mem[9898] = 126;
razn_h_mem[9899] = 2;
razn_h_mem[9900] = 132;
razn_h_mem[9901] = 8;
razn_h_mem[9902] = 138;
razn_h_mem[9903] = 14;
razn_h_mem[9904] = 144;
razn_h_mem[9905] = 20;
razn_h_mem[9906] = 150;
razn_h_mem[9907] = 26;
razn_h_mem[9908] = 156;
razn_h_mem[9909] = 32;
razn_h_mem[9910] = 162;
razn_h_mem[9911] = 38;
razn_h_mem[9912] = 168;
razn_h_mem[9913] = 44;
razn_h_mem[9914] = 174;
razn_h_mem[9915] = 50;
razn_h_mem[9916] = 180;
razn_h_mem[9917] = 56;
razn_h_mem[9918] = 186;
razn_h_mem[9919] = 62;
razn_h_mem[9920] = 192;
razn_h_mem[9921] = 68;
razn_h_mem[9922] = 198;
razn_h_mem[9923] = 74;
razn_h_mem[9924] = 204;
razn_h_mem[9925] = 80;
razn_h_mem[9926] = 210;
razn_h_mem[9927] = 86;
razn_h_mem[9928] = 216;
razn_h_mem[9929] = 92;
razn_h_mem[9930] = 222;
razn_h_mem[9931] = 98;
razn_h_mem[9932] = 228;
razn_h_mem[9933] = 104;
razn_h_mem[9934] = 234;
razn_h_mem[9935] = 110;
razn_h_mem[9936] = 240;
razn_h_mem[9937] = 116;
razn_h_mem[9938] = 246;
razn_h_mem[9939] = 122;
razn_h_mem[9940] = 252;
razn_h_mem[9941] = 128;
razn_h_mem[9942] = 4;
razn_h_mem[9943] = 134;
razn_h_mem[9944] = 10;
razn_h_mem[9945] = 140;
razn_h_mem[9946] = 16;
razn_h_mem[9947] = 146;
razn_h_mem[9948] = 22;
razn_h_mem[9949] = 152;
razn_h_mem[9950] = 28;
razn_h_mem[9951] = 158;
razn_h_mem[9952] = 34;
razn_h_mem[9953] = 164;
razn_h_mem[9954] = 40;
razn_h_mem[9955] = 170;
razn_h_mem[9956] = 46;
razn_h_mem[9957] = 176;
razn_h_mem[9958] = 52;
razn_h_mem[9959] = 182;
razn_h_mem[9960] = 58;
razn_h_mem[9961] = 188;
razn_h_mem[9962] = 64;
razn_h_mem[9963] = 194;
razn_h_mem[9964] = 70;
razn_h_mem[9965] = 200;
razn_h_mem[9966] = 76;
razn_h_mem[9967] = 206;
razn_h_mem[9968] = 82;
razn_h_mem[9969] = 212;
razn_h_mem[9970] = 88;
razn_h_mem[9971] = 218;
razn_h_mem[9972] = 94;
razn_h_mem[9973] = 224;
razn_h_mem[9974] = 100;
razn_h_mem[9975] = 230;
razn_h_mem[9976] = 106;
razn_h_mem[9977] = 236;
razn_h_mem[9978] = 112;
razn_h_mem[9979] = 242;
razn_h_mem[9980] = 118;
razn_h_mem[9981] = 248;
razn_h_mem[9982] = 124;
razn_h_mem[9983] = 255;
razn_h_mem[9984] = 0;
razn_h_mem[9985] = 130;
razn_h_mem[9986] = 6;
razn_h_mem[9987] = 136;
razn_h_mem[9988] = 12;
razn_h_mem[9989] = 142;
razn_h_mem[9990] = 18;
razn_h_mem[9991] = 148;
razn_h_mem[9992] = 24;
razn_h_mem[9993] = 154;
razn_h_mem[9994] = 30;
razn_h_mem[9995] = 160;
razn_h_mem[9996] = 36;
razn_h_mem[9997] = 166;
razn_h_mem[9998] = 42;
razn_h_mem[9999] = 172;
razn_h_mem[10000] = 48;
razn_h_mem[10001] = 178;
razn_h_mem[10002] = 54;
razn_h_mem[10003] = 184;
razn_h_mem[10004] = 60;
razn_h_mem[10005] = 190;
razn_h_mem[10006] = 66;
razn_h_mem[10007] = 196;
razn_h_mem[10008] = 72;
razn_h_mem[10009] = 202;
razn_h_mem[10010] = 78;
razn_h_mem[10011] = 208;
razn_h_mem[10012] = 84;
razn_h_mem[10013] = 214;
razn_h_mem[10014] = 90;
razn_h_mem[10015] = 220;
razn_h_mem[10016] = 96;
razn_h_mem[10017] = 226;
razn_h_mem[10018] = 102;
razn_h_mem[10019] = 232;
razn_h_mem[10020] = 108;
razn_h_mem[10021] = 238;
razn_h_mem[10022] = 114;
razn_h_mem[10023] = 244;
razn_h_mem[10024] = 120;
razn_h_mem[10025] = 250;
razn_h_mem[10026] = 126;
razn_h_mem[10027] = 2;
razn_h_mem[10028] = 132;
razn_h_mem[10029] = 8;
razn_h_mem[10030] = 138;
razn_h_mem[10031] = 14;
razn_h_mem[10032] = 144;
razn_h_mem[10033] = 20;
razn_h_mem[10034] = 150;
razn_h_mem[10035] = 26;
razn_h_mem[10036] = 156;
razn_h_mem[10037] = 32;
razn_h_mem[10038] = 162;
razn_h_mem[10039] = 38;
razn_h_mem[10040] = 168;
razn_h_mem[10041] = 44;
razn_h_mem[10042] = 174;
razn_h_mem[10043] = 50;
razn_h_mem[10044] = 180;
razn_h_mem[10045] = 56;
razn_h_mem[10046] = 186;
razn_h_mem[10047] = 62;
razn_h_mem[10048] = 192;
razn_h_mem[10049] = 68;
razn_h_mem[10050] = 198;
razn_h_mem[10051] = 74;
razn_h_mem[10052] = 204;
razn_h_mem[10053] = 80;
razn_h_mem[10054] = 210;
razn_h_mem[10055] = 86;
razn_h_mem[10056] = 216;
razn_h_mem[10057] = 92;
razn_h_mem[10058] = 222;
razn_h_mem[10059] = 98;
razn_h_mem[10060] = 228;
razn_h_mem[10061] = 104;
razn_h_mem[10062] = 234;
razn_h_mem[10063] = 110;
razn_h_mem[10064] = 240;
razn_h_mem[10065] = 116;
razn_h_mem[10066] = 246;
razn_h_mem[10067] = 122;
razn_h_mem[10068] = 252;
razn_h_mem[10069] = 128;
razn_h_mem[10070] = 4;
razn_h_mem[10071] = 134;
razn_h_mem[10072] = 10;
razn_h_mem[10073] = 140;
razn_h_mem[10074] = 16;
razn_h_mem[10075] = 146;
razn_h_mem[10076] = 22;
razn_h_mem[10077] = 152;
razn_h_mem[10078] = 28;
razn_h_mem[10079] = 158;
razn_h_mem[10080] = 34;
razn_h_mem[10081] = 164;
razn_h_mem[10082] = 40;
razn_h_mem[10083] = 170;
razn_h_mem[10084] = 46;
razn_h_mem[10085] = 176;
razn_h_mem[10086] = 52;
razn_h_mem[10087] = 182;
razn_h_mem[10088] = 58;
razn_h_mem[10089] = 188;
razn_h_mem[10090] = 64;
razn_h_mem[10091] = 194;
razn_h_mem[10092] = 70;
razn_h_mem[10093] = 200;
razn_h_mem[10094] = 76;
razn_h_mem[10095] = 206;
razn_h_mem[10096] = 82;
razn_h_mem[10097] = 212;
razn_h_mem[10098] = 88;
razn_h_mem[10099] = 218;
razn_h_mem[10100] = 94;
razn_h_mem[10101] = 224;
razn_h_mem[10102] = 100;
razn_h_mem[10103] = 230;
razn_h_mem[10104] = 106;
razn_h_mem[10105] = 236;
razn_h_mem[10106] = 112;
razn_h_mem[10107] = 242;
razn_h_mem[10108] = 118;
razn_h_mem[10109] = 248;
razn_h_mem[10110] = 124;
razn_h_mem[10111] = 255;
razn_h_mem[10112] = 0;
razn_h_mem[10113] = 130;
razn_h_mem[10114] = 6;
razn_h_mem[10115] = 136;
razn_h_mem[10116] = 12;
razn_h_mem[10117] = 142;
razn_h_mem[10118] = 18;
razn_h_mem[10119] = 148;
razn_h_mem[10120] = 24;
razn_h_mem[10121] = 154;
razn_h_mem[10122] = 30;
razn_h_mem[10123] = 160;
razn_h_mem[10124] = 36;
razn_h_mem[10125] = 166;
razn_h_mem[10126] = 42;
razn_h_mem[10127] = 172;
razn_h_mem[10128] = 48;
razn_h_mem[10129] = 178;
razn_h_mem[10130] = 54;
razn_h_mem[10131] = 184;
razn_h_mem[10132] = 60;
razn_h_mem[10133] = 190;
razn_h_mem[10134] = 66;
razn_h_mem[10135] = 196;
razn_h_mem[10136] = 72;
razn_h_mem[10137] = 202;
razn_h_mem[10138] = 78;
razn_h_mem[10139] = 208;
razn_h_mem[10140] = 84;
razn_h_mem[10141] = 214;
razn_h_mem[10142] = 90;
razn_h_mem[10143] = 220;
razn_h_mem[10144] = 96;
razn_h_mem[10145] = 226;
razn_h_mem[10146] = 102;
razn_h_mem[10147] = 232;
razn_h_mem[10148] = 108;
razn_h_mem[10149] = 238;
razn_h_mem[10150] = 114;
razn_h_mem[10151] = 244;
razn_h_mem[10152] = 120;
razn_h_mem[10153] = 250;
razn_h_mem[10154] = 126;
razn_h_mem[10155] = 2;
razn_h_mem[10156] = 132;
razn_h_mem[10157] = 8;
razn_h_mem[10158] = 138;
razn_h_mem[10159] = 14;
razn_h_mem[10160] = 144;
razn_h_mem[10161] = 20;
razn_h_mem[10162] = 150;
razn_h_mem[10163] = 26;
razn_h_mem[10164] = 156;
razn_h_mem[10165] = 32;
razn_h_mem[10166] = 162;
razn_h_mem[10167] = 38;
razn_h_mem[10168] = 168;
razn_h_mem[10169] = 44;
razn_h_mem[10170] = 174;
razn_h_mem[10171] = 50;
razn_h_mem[10172] = 180;
razn_h_mem[10173] = 56;
razn_h_mem[10174] = 186;
razn_h_mem[10175] = 62;
razn_h_mem[10176] = 192;
razn_h_mem[10177] = 68;
razn_h_mem[10178] = 198;
razn_h_mem[10179] = 74;
razn_h_mem[10180] = 204;
razn_h_mem[10181] = 80;
razn_h_mem[10182] = 210;
razn_h_mem[10183] = 86;
razn_h_mem[10184] = 216;
razn_h_mem[10185] = 92;
razn_h_mem[10186] = 222;
razn_h_mem[10187] = 98;
razn_h_mem[10188] = 228;
razn_h_mem[10189] = 104;
razn_h_mem[10190] = 234;
razn_h_mem[10191] = 110;
razn_h_mem[10192] = 240;
razn_h_mem[10193] = 116;
razn_h_mem[10194] = 246;
razn_h_mem[10195] = 122;
razn_h_mem[10196] = 252;
razn_h_mem[10197] = 128;
razn_h_mem[10198] = 4;
razn_h_mem[10199] = 134;
razn_h_mem[10200] = 10;
razn_h_mem[10201] = 140;
razn_h_mem[10202] = 16;
razn_h_mem[10203] = 146;
razn_h_mem[10204] = 22;
razn_h_mem[10205] = 152;
razn_h_mem[10206] = 28;
razn_h_mem[10207] = 158;
razn_h_mem[10208] = 34;
razn_h_mem[10209] = 164;
razn_h_mem[10210] = 40;
razn_h_mem[10211] = 170;
razn_h_mem[10212] = 46;
razn_h_mem[10213] = 176;
razn_h_mem[10214] = 52;
razn_h_mem[10215] = 182;
razn_h_mem[10216] = 58;
razn_h_mem[10217] = 188;
razn_h_mem[10218] = 64;
razn_h_mem[10219] = 194;
razn_h_mem[10220] = 70;
razn_h_mem[10221] = 200;
razn_h_mem[10222] = 76;
razn_h_mem[10223] = 206;
razn_h_mem[10224] = 82;
razn_h_mem[10225] = 212;
razn_h_mem[10226] = 88;
razn_h_mem[10227] = 218;
razn_h_mem[10228] = 94;
razn_h_mem[10229] = 224;
razn_h_mem[10230] = 100;
razn_h_mem[10231] = 230;
razn_h_mem[10232] = 106;
razn_h_mem[10233] = 236;
razn_h_mem[10234] = 112;
razn_h_mem[10235] = 242;
razn_h_mem[10236] = 118;
razn_h_mem[10237] = 248;
razn_h_mem[10238] = 124;
razn_h_mem[10239] = 255;
razn_h_mem[10240] = 0;
razn_h_mem[10241] = 130;
razn_h_mem[10242] = 6;
razn_h_mem[10243] = 136;
razn_h_mem[10244] = 12;
razn_h_mem[10245] = 142;
razn_h_mem[10246] = 18;
razn_h_mem[10247] = 148;
razn_h_mem[10248] = 24;
razn_h_mem[10249] = 154;
razn_h_mem[10250] = 30;
razn_h_mem[10251] = 160;
razn_h_mem[10252] = 36;
razn_h_mem[10253] = 166;
razn_h_mem[10254] = 42;
razn_h_mem[10255] = 172;
razn_h_mem[10256] = 48;
razn_h_mem[10257] = 178;
razn_h_mem[10258] = 54;
razn_h_mem[10259] = 184;
razn_h_mem[10260] = 60;
razn_h_mem[10261] = 190;
razn_h_mem[10262] = 66;
razn_h_mem[10263] = 196;
razn_h_mem[10264] = 72;
razn_h_mem[10265] = 202;
razn_h_mem[10266] = 78;
razn_h_mem[10267] = 208;
razn_h_mem[10268] = 84;
razn_h_mem[10269] = 214;
razn_h_mem[10270] = 90;
razn_h_mem[10271] = 220;
razn_h_mem[10272] = 96;
razn_h_mem[10273] = 226;
razn_h_mem[10274] = 102;
razn_h_mem[10275] = 232;
razn_h_mem[10276] = 108;
razn_h_mem[10277] = 238;
razn_h_mem[10278] = 114;
razn_h_mem[10279] = 244;
razn_h_mem[10280] = 120;
razn_h_mem[10281] = 250;
razn_h_mem[10282] = 126;
razn_h_mem[10283] = 2;
razn_h_mem[10284] = 132;
razn_h_mem[10285] = 8;
razn_h_mem[10286] = 138;
razn_h_mem[10287] = 14;
razn_h_mem[10288] = 144;
razn_h_mem[10289] = 20;
razn_h_mem[10290] = 150;
razn_h_mem[10291] = 26;
razn_h_mem[10292] = 156;
razn_h_mem[10293] = 32;
razn_h_mem[10294] = 162;
razn_h_mem[10295] = 38;
razn_h_mem[10296] = 168;
razn_h_mem[10297] = 44;
razn_h_mem[10298] = 174;
razn_h_mem[10299] = 50;
razn_h_mem[10300] = 180;
razn_h_mem[10301] = 56;
razn_h_mem[10302] = 186;
razn_h_mem[10303] = 62;
razn_h_mem[10304] = 192;
razn_h_mem[10305] = 68;
razn_h_mem[10306] = 198;
razn_h_mem[10307] = 74;
razn_h_mem[10308] = 204;
razn_h_mem[10309] = 80;
razn_h_mem[10310] = 210;
razn_h_mem[10311] = 86;
razn_h_mem[10312] = 216;
razn_h_mem[10313] = 92;
razn_h_mem[10314] = 222;
razn_h_mem[10315] = 98;
razn_h_mem[10316] = 228;
razn_h_mem[10317] = 104;
razn_h_mem[10318] = 234;
razn_h_mem[10319] = 110;
razn_h_mem[10320] = 240;
razn_h_mem[10321] = 116;
razn_h_mem[10322] = 246;
razn_h_mem[10323] = 122;
razn_h_mem[10324] = 252;
razn_h_mem[10325] = 128;
razn_h_mem[10326] = 4;
razn_h_mem[10327] = 134;
razn_h_mem[10328] = 10;
razn_h_mem[10329] = 140;
razn_h_mem[10330] = 16;
razn_h_mem[10331] = 146;
razn_h_mem[10332] = 22;
razn_h_mem[10333] = 152;
razn_h_mem[10334] = 28;
razn_h_mem[10335] = 158;
razn_h_mem[10336] = 34;
razn_h_mem[10337] = 164;
razn_h_mem[10338] = 40;
razn_h_mem[10339] = 170;
razn_h_mem[10340] = 46;
razn_h_mem[10341] = 176;
razn_h_mem[10342] = 52;
razn_h_mem[10343] = 182;
razn_h_mem[10344] = 58;
razn_h_mem[10345] = 188;
razn_h_mem[10346] = 64;
razn_h_mem[10347] = 194;
razn_h_mem[10348] = 70;
razn_h_mem[10349] = 200;
razn_h_mem[10350] = 76;
razn_h_mem[10351] = 206;
razn_h_mem[10352] = 82;
razn_h_mem[10353] = 212;
razn_h_mem[10354] = 88;
razn_h_mem[10355] = 218;
razn_h_mem[10356] = 94;
razn_h_mem[10357] = 224;
razn_h_mem[10358] = 100;
razn_h_mem[10359] = 230;
razn_h_mem[10360] = 106;
razn_h_mem[10361] = 236;
razn_h_mem[10362] = 112;
razn_h_mem[10363] = 242;
razn_h_mem[10364] = 118;
razn_h_mem[10365] = 248;
razn_h_mem[10366] = 124;
razn_h_mem[10367] = 255;
razn_h_mem[10368] = 0;
razn_h_mem[10369] = 130;
razn_h_mem[10370] = 6;
razn_h_mem[10371] = 136;
razn_h_mem[10372] = 12;
razn_h_mem[10373] = 142;
razn_h_mem[10374] = 18;
razn_h_mem[10375] = 148;
razn_h_mem[10376] = 24;
razn_h_mem[10377] = 154;
razn_h_mem[10378] = 30;
razn_h_mem[10379] = 160;
razn_h_mem[10380] = 36;
razn_h_mem[10381] = 166;
razn_h_mem[10382] = 42;
razn_h_mem[10383] = 172;
razn_h_mem[10384] = 48;
razn_h_mem[10385] = 178;
razn_h_mem[10386] = 54;
razn_h_mem[10387] = 184;
razn_h_mem[10388] = 60;
razn_h_mem[10389] = 190;
razn_h_mem[10390] = 66;
razn_h_mem[10391] = 196;
razn_h_mem[10392] = 72;
razn_h_mem[10393] = 202;
razn_h_mem[10394] = 78;
razn_h_mem[10395] = 208;
razn_h_mem[10396] = 84;
razn_h_mem[10397] = 214;
razn_h_mem[10398] = 90;
razn_h_mem[10399] = 220;
razn_h_mem[10400] = 96;
razn_h_mem[10401] = 226;
razn_h_mem[10402] = 102;
razn_h_mem[10403] = 232;
razn_h_mem[10404] = 108;
razn_h_mem[10405] = 238;
razn_h_mem[10406] = 114;
razn_h_mem[10407] = 244;
razn_h_mem[10408] = 120;
razn_h_mem[10409] = 250;
razn_h_mem[10410] = 126;
razn_h_mem[10411] = 2;
razn_h_mem[10412] = 132;
razn_h_mem[10413] = 8;
razn_h_mem[10414] = 138;
razn_h_mem[10415] = 14;
razn_h_mem[10416] = 144;
razn_h_mem[10417] = 20;
razn_h_mem[10418] = 150;
razn_h_mem[10419] = 26;
razn_h_mem[10420] = 156;
razn_h_mem[10421] = 32;
razn_h_mem[10422] = 162;
razn_h_mem[10423] = 38;
razn_h_mem[10424] = 168;
razn_h_mem[10425] = 44;
razn_h_mem[10426] = 174;
razn_h_mem[10427] = 50;
razn_h_mem[10428] = 180;
razn_h_mem[10429] = 56;
razn_h_mem[10430] = 186;
razn_h_mem[10431] = 62;
razn_h_mem[10432] = 192;
razn_h_mem[10433] = 68;
razn_h_mem[10434] = 198;
razn_h_mem[10435] = 74;
razn_h_mem[10436] = 204;
razn_h_mem[10437] = 80;
razn_h_mem[10438] = 210;
razn_h_mem[10439] = 86;
razn_h_mem[10440] = 216;
razn_h_mem[10441] = 92;
razn_h_mem[10442] = 222;
razn_h_mem[10443] = 98;
razn_h_mem[10444] = 228;
razn_h_mem[10445] = 104;
razn_h_mem[10446] = 234;
razn_h_mem[10447] = 110;
razn_h_mem[10448] = 240;
razn_h_mem[10449] = 116;
razn_h_mem[10450] = 246;
razn_h_mem[10451] = 122;
razn_h_mem[10452] = 252;
razn_h_mem[10453] = 128;
razn_h_mem[10454] = 4;
razn_h_mem[10455] = 134;
razn_h_mem[10456] = 10;
razn_h_mem[10457] = 140;
razn_h_mem[10458] = 16;
razn_h_mem[10459] = 146;
razn_h_mem[10460] = 22;
razn_h_mem[10461] = 152;
razn_h_mem[10462] = 28;
razn_h_mem[10463] = 158;
razn_h_mem[10464] = 34;
razn_h_mem[10465] = 164;
razn_h_mem[10466] = 40;
razn_h_mem[10467] = 170;
razn_h_mem[10468] = 46;
razn_h_mem[10469] = 176;
razn_h_mem[10470] = 52;
razn_h_mem[10471] = 182;
razn_h_mem[10472] = 58;
razn_h_mem[10473] = 188;
razn_h_mem[10474] = 64;
razn_h_mem[10475] = 194;
razn_h_mem[10476] = 70;
razn_h_mem[10477] = 200;
razn_h_mem[10478] = 76;
razn_h_mem[10479] = 206;
razn_h_mem[10480] = 82;
razn_h_mem[10481] = 212;
razn_h_mem[10482] = 88;
razn_h_mem[10483] = 218;
razn_h_mem[10484] = 94;
razn_h_mem[10485] = 224;
razn_h_mem[10486] = 100;
razn_h_mem[10487] = 230;
razn_h_mem[10488] = 106;
razn_h_mem[10489] = 236;
razn_h_mem[10490] = 112;
razn_h_mem[10491] = 242;
razn_h_mem[10492] = 118;
razn_h_mem[10493] = 248;
razn_h_mem[10494] = 124;
razn_h_mem[10495] = 255;
razn_h_mem[10496] = 0;
razn_h_mem[10497] = 130;
razn_h_mem[10498] = 6;
razn_h_mem[10499] = 136;
razn_h_mem[10500] = 12;
razn_h_mem[10501] = 142;
razn_h_mem[10502] = 18;
razn_h_mem[10503] = 148;
razn_h_mem[10504] = 24;
razn_h_mem[10505] = 154;
razn_h_mem[10506] = 30;
razn_h_mem[10507] = 160;
razn_h_mem[10508] = 36;
razn_h_mem[10509] = 166;
razn_h_mem[10510] = 42;
razn_h_mem[10511] = 172;
razn_h_mem[10512] = 48;
razn_h_mem[10513] = 178;
razn_h_mem[10514] = 54;
razn_h_mem[10515] = 184;
razn_h_mem[10516] = 60;
razn_h_mem[10517] = 190;
razn_h_mem[10518] = 66;
razn_h_mem[10519] = 196;
razn_h_mem[10520] = 72;
razn_h_mem[10521] = 202;
razn_h_mem[10522] = 78;
razn_h_mem[10523] = 208;
razn_h_mem[10524] = 84;
razn_h_mem[10525] = 214;
razn_h_mem[10526] = 90;
razn_h_mem[10527] = 220;
razn_h_mem[10528] = 96;
razn_h_mem[10529] = 226;
razn_h_mem[10530] = 102;
razn_h_mem[10531] = 232;
razn_h_mem[10532] = 108;
razn_h_mem[10533] = 238;
razn_h_mem[10534] = 114;
razn_h_mem[10535] = 244;
razn_h_mem[10536] = 120;
razn_h_mem[10537] = 250;
razn_h_mem[10538] = 126;
razn_h_mem[10539] = 2;
razn_h_mem[10540] = 132;
razn_h_mem[10541] = 8;
razn_h_mem[10542] = 138;
razn_h_mem[10543] = 14;
razn_h_mem[10544] = 144;
razn_h_mem[10545] = 20;
razn_h_mem[10546] = 150;
razn_h_mem[10547] = 26;
razn_h_mem[10548] = 156;
razn_h_mem[10549] = 32;
razn_h_mem[10550] = 162;
razn_h_mem[10551] = 38;
razn_h_mem[10552] = 168;
razn_h_mem[10553] = 44;
razn_h_mem[10554] = 174;
razn_h_mem[10555] = 50;
razn_h_mem[10556] = 180;
razn_h_mem[10557] = 56;
razn_h_mem[10558] = 186;
razn_h_mem[10559] = 62;
razn_h_mem[10560] = 192;
razn_h_mem[10561] = 68;
razn_h_mem[10562] = 198;
razn_h_mem[10563] = 74;
razn_h_mem[10564] = 204;
razn_h_mem[10565] = 80;
razn_h_mem[10566] = 210;
razn_h_mem[10567] = 86;
razn_h_mem[10568] = 216;
razn_h_mem[10569] = 92;
razn_h_mem[10570] = 222;
razn_h_mem[10571] = 98;
razn_h_mem[10572] = 228;
razn_h_mem[10573] = 104;
razn_h_mem[10574] = 234;
razn_h_mem[10575] = 110;
razn_h_mem[10576] = 240;
razn_h_mem[10577] = 116;
razn_h_mem[10578] = 246;
razn_h_mem[10579] = 122;
razn_h_mem[10580] = 252;
razn_h_mem[10581] = 128;
razn_h_mem[10582] = 4;
razn_h_mem[10583] = 134;
razn_h_mem[10584] = 10;
razn_h_mem[10585] = 140;
razn_h_mem[10586] = 16;
razn_h_mem[10587] = 146;
razn_h_mem[10588] = 22;
razn_h_mem[10589] = 152;
razn_h_mem[10590] = 28;
razn_h_mem[10591] = 158;
razn_h_mem[10592] = 34;
razn_h_mem[10593] = 164;
razn_h_mem[10594] = 40;
razn_h_mem[10595] = 170;
razn_h_mem[10596] = 46;
razn_h_mem[10597] = 176;
razn_h_mem[10598] = 52;
razn_h_mem[10599] = 182;
razn_h_mem[10600] = 58;
razn_h_mem[10601] = 188;
razn_h_mem[10602] = 64;
razn_h_mem[10603] = 194;
razn_h_mem[10604] = 70;
razn_h_mem[10605] = 200;
razn_h_mem[10606] = 76;
razn_h_mem[10607] = 206;
razn_h_mem[10608] = 82;
razn_h_mem[10609] = 212;
razn_h_mem[10610] = 88;
razn_h_mem[10611] = 218;
razn_h_mem[10612] = 94;
razn_h_mem[10613] = 224;
razn_h_mem[10614] = 100;
razn_h_mem[10615] = 230;
razn_h_mem[10616] = 106;
razn_h_mem[10617] = 236;
razn_h_mem[10618] = 112;
razn_h_mem[10619] = 242;
razn_h_mem[10620] = 118;
razn_h_mem[10621] = 248;
razn_h_mem[10622] = 124;
razn_h_mem[10623] = 255;
razn_h_mem[10624] = 0;
razn_h_mem[10625] = 130;
razn_h_mem[10626] = 6;
razn_h_mem[10627] = 136;
razn_h_mem[10628] = 12;
razn_h_mem[10629] = 142;
razn_h_mem[10630] = 18;
razn_h_mem[10631] = 148;
razn_h_mem[10632] = 24;
razn_h_mem[10633] = 154;
razn_h_mem[10634] = 30;
razn_h_mem[10635] = 160;
razn_h_mem[10636] = 36;
razn_h_mem[10637] = 166;
razn_h_mem[10638] = 42;
razn_h_mem[10639] = 172;
razn_h_mem[10640] = 48;
razn_h_mem[10641] = 178;
razn_h_mem[10642] = 54;
razn_h_mem[10643] = 184;
razn_h_mem[10644] = 60;
razn_h_mem[10645] = 190;
razn_h_mem[10646] = 66;
razn_h_mem[10647] = 196;
razn_h_mem[10648] = 72;
razn_h_mem[10649] = 202;
razn_h_mem[10650] = 78;
razn_h_mem[10651] = 208;
razn_h_mem[10652] = 84;
razn_h_mem[10653] = 214;
razn_h_mem[10654] = 90;
razn_h_mem[10655] = 220;
razn_h_mem[10656] = 96;
razn_h_mem[10657] = 226;
razn_h_mem[10658] = 102;
razn_h_mem[10659] = 232;
razn_h_mem[10660] = 108;
razn_h_mem[10661] = 238;
razn_h_mem[10662] = 114;
razn_h_mem[10663] = 244;
razn_h_mem[10664] = 120;
razn_h_mem[10665] = 250;
razn_h_mem[10666] = 126;
razn_h_mem[10667] = 2;
razn_h_mem[10668] = 132;
razn_h_mem[10669] = 8;
razn_h_mem[10670] = 138;
razn_h_mem[10671] = 14;
razn_h_mem[10672] = 144;
razn_h_mem[10673] = 20;
razn_h_mem[10674] = 150;
razn_h_mem[10675] = 26;
razn_h_mem[10676] = 156;
razn_h_mem[10677] = 32;
razn_h_mem[10678] = 162;
razn_h_mem[10679] = 38;
razn_h_mem[10680] = 168;
razn_h_mem[10681] = 44;
razn_h_mem[10682] = 174;
razn_h_mem[10683] = 50;
razn_h_mem[10684] = 180;
razn_h_mem[10685] = 56;
razn_h_mem[10686] = 186;
razn_h_mem[10687] = 62;
razn_h_mem[10688] = 192;
razn_h_mem[10689] = 68;
razn_h_mem[10690] = 198;
razn_h_mem[10691] = 74;
razn_h_mem[10692] = 204;
razn_h_mem[10693] = 80;
razn_h_mem[10694] = 210;
razn_h_mem[10695] = 86;
razn_h_mem[10696] = 216;
razn_h_mem[10697] = 92;
razn_h_mem[10698] = 222;
razn_h_mem[10699] = 98;
razn_h_mem[10700] = 228;
razn_h_mem[10701] = 104;
razn_h_mem[10702] = 234;
razn_h_mem[10703] = 110;
razn_h_mem[10704] = 240;
razn_h_mem[10705] = 116;
razn_h_mem[10706] = 246;
razn_h_mem[10707] = 122;
razn_h_mem[10708] = 252;
razn_h_mem[10709] = 128;
razn_h_mem[10710] = 4;
razn_h_mem[10711] = 134;
razn_h_mem[10712] = 10;
razn_h_mem[10713] = 140;
razn_h_mem[10714] = 16;
razn_h_mem[10715] = 146;
razn_h_mem[10716] = 22;
razn_h_mem[10717] = 152;
razn_h_mem[10718] = 28;
razn_h_mem[10719] = 158;
razn_h_mem[10720] = 34;
razn_h_mem[10721] = 164;
razn_h_mem[10722] = 40;
razn_h_mem[10723] = 170;
razn_h_mem[10724] = 46;
razn_h_mem[10725] = 176;
razn_h_mem[10726] = 52;
razn_h_mem[10727] = 182;
razn_h_mem[10728] = 58;
razn_h_mem[10729] = 188;
razn_h_mem[10730] = 64;
razn_h_mem[10731] = 194;
razn_h_mem[10732] = 70;
razn_h_mem[10733] = 200;
razn_h_mem[10734] = 76;
razn_h_mem[10735] = 206;
razn_h_mem[10736] = 82;
razn_h_mem[10737] = 212;
razn_h_mem[10738] = 88;
razn_h_mem[10739] = 218;
razn_h_mem[10740] = 94;
razn_h_mem[10741] = 224;
razn_h_mem[10742] = 100;
razn_h_mem[10743] = 230;
razn_h_mem[10744] = 106;
razn_h_mem[10745] = 236;
razn_h_mem[10746] = 112;
razn_h_mem[10747] = 242;
razn_h_mem[10748] = 118;
razn_h_mem[10749] = 248;
razn_h_mem[10750] = 124;
razn_h_mem[10751] = 255;
razn_h_mem[10752] = 0;
razn_h_mem[10753] = 130;
razn_h_mem[10754] = 6;
razn_h_mem[10755] = 136;
razn_h_mem[10756] = 12;
razn_h_mem[10757] = 142;
razn_h_mem[10758] = 18;
razn_h_mem[10759] = 148;
razn_h_mem[10760] = 24;
razn_h_mem[10761] = 154;
razn_h_mem[10762] = 30;
razn_h_mem[10763] = 160;
razn_h_mem[10764] = 36;
razn_h_mem[10765] = 166;
razn_h_mem[10766] = 42;
razn_h_mem[10767] = 172;
razn_h_mem[10768] = 48;
razn_h_mem[10769] = 178;
razn_h_mem[10770] = 54;
razn_h_mem[10771] = 184;
razn_h_mem[10772] = 60;
razn_h_mem[10773] = 190;
razn_h_mem[10774] = 66;
razn_h_mem[10775] = 196;
razn_h_mem[10776] = 72;
razn_h_mem[10777] = 202;
razn_h_mem[10778] = 78;
razn_h_mem[10779] = 208;
razn_h_mem[10780] = 84;
razn_h_mem[10781] = 214;
razn_h_mem[10782] = 90;
razn_h_mem[10783] = 220;
razn_h_mem[10784] = 96;
razn_h_mem[10785] = 226;
razn_h_mem[10786] = 102;
razn_h_mem[10787] = 232;
razn_h_mem[10788] = 108;
razn_h_mem[10789] = 238;
razn_h_mem[10790] = 114;
razn_h_mem[10791] = 244;
razn_h_mem[10792] = 120;
razn_h_mem[10793] = 250;
razn_h_mem[10794] = 126;
razn_h_mem[10795] = 2;
razn_h_mem[10796] = 132;
razn_h_mem[10797] = 8;
razn_h_mem[10798] = 138;
razn_h_mem[10799] = 14;
razn_h_mem[10800] = 144;
razn_h_mem[10801] = 20;
razn_h_mem[10802] = 150;
razn_h_mem[10803] = 26;
razn_h_mem[10804] = 156;
razn_h_mem[10805] = 32;
razn_h_mem[10806] = 162;
razn_h_mem[10807] = 38;
razn_h_mem[10808] = 168;
razn_h_mem[10809] = 44;
razn_h_mem[10810] = 174;
razn_h_mem[10811] = 50;
razn_h_mem[10812] = 180;
razn_h_mem[10813] = 56;
razn_h_mem[10814] = 186;
razn_h_mem[10815] = 62;
razn_h_mem[10816] = 192;
razn_h_mem[10817] = 68;
razn_h_mem[10818] = 198;
razn_h_mem[10819] = 74;
razn_h_mem[10820] = 204;
razn_h_mem[10821] = 80;
razn_h_mem[10822] = 210;
razn_h_mem[10823] = 86;
razn_h_mem[10824] = 216;
razn_h_mem[10825] = 92;
razn_h_mem[10826] = 222;
razn_h_mem[10827] = 98;
razn_h_mem[10828] = 228;
razn_h_mem[10829] = 104;
razn_h_mem[10830] = 234;
razn_h_mem[10831] = 110;
razn_h_mem[10832] = 240;
razn_h_mem[10833] = 116;
razn_h_mem[10834] = 246;
razn_h_mem[10835] = 122;
razn_h_mem[10836] = 252;
razn_h_mem[10837] = 128;
razn_h_mem[10838] = 4;
razn_h_mem[10839] = 134;
razn_h_mem[10840] = 10;
razn_h_mem[10841] = 140;
razn_h_mem[10842] = 16;
razn_h_mem[10843] = 146;
razn_h_mem[10844] = 22;
razn_h_mem[10845] = 152;
razn_h_mem[10846] = 28;
razn_h_mem[10847] = 158;
razn_h_mem[10848] = 34;
razn_h_mem[10849] = 164;
razn_h_mem[10850] = 40;
razn_h_mem[10851] = 170;
razn_h_mem[10852] = 46;
razn_h_mem[10853] = 176;
razn_h_mem[10854] = 52;
razn_h_mem[10855] = 182;
razn_h_mem[10856] = 58;
razn_h_mem[10857] = 188;
razn_h_mem[10858] = 64;
razn_h_mem[10859] = 194;
razn_h_mem[10860] = 70;
razn_h_mem[10861] = 200;
razn_h_mem[10862] = 76;
razn_h_mem[10863] = 206;
razn_h_mem[10864] = 82;
razn_h_mem[10865] = 212;
razn_h_mem[10866] = 88;
razn_h_mem[10867] = 218;
razn_h_mem[10868] = 94;
razn_h_mem[10869] = 224;
razn_h_mem[10870] = 100;
razn_h_mem[10871] = 230;
razn_h_mem[10872] = 106;
razn_h_mem[10873] = 236;
razn_h_mem[10874] = 112;
razn_h_mem[10875] = 242;
razn_h_mem[10876] = 118;
razn_h_mem[10877] = 248;
razn_h_mem[10878] = 124;
razn_h_mem[10879] = 255;
razn_h_mem[10880] = 0;
razn_h_mem[10881] = 130;
razn_h_mem[10882] = 6;
razn_h_mem[10883] = 136;
razn_h_mem[10884] = 12;
razn_h_mem[10885] = 142;
razn_h_mem[10886] = 18;
razn_h_mem[10887] = 148;
razn_h_mem[10888] = 24;
razn_h_mem[10889] = 154;
razn_h_mem[10890] = 30;
razn_h_mem[10891] = 160;
razn_h_mem[10892] = 36;
razn_h_mem[10893] = 166;
razn_h_mem[10894] = 42;
razn_h_mem[10895] = 172;
razn_h_mem[10896] = 48;
razn_h_mem[10897] = 178;
razn_h_mem[10898] = 54;
razn_h_mem[10899] = 184;
razn_h_mem[10900] = 60;
razn_h_mem[10901] = 190;
razn_h_mem[10902] = 66;
razn_h_mem[10903] = 196;
razn_h_mem[10904] = 72;
razn_h_mem[10905] = 202;
razn_h_mem[10906] = 78;
razn_h_mem[10907] = 208;
razn_h_mem[10908] = 84;
razn_h_mem[10909] = 214;
razn_h_mem[10910] = 90;
razn_h_mem[10911] = 220;
razn_h_mem[10912] = 96;
razn_h_mem[10913] = 226;
razn_h_mem[10914] = 102;
razn_h_mem[10915] = 232;
razn_h_mem[10916] = 108;
razn_h_mem[10917] = 238;
razn_h_mem[10918] = 114;
razn_h_mem[10919] = 244;
razn_h_mem[10920] = 120;
razn_h_mem[10921] = 250;
razn_h_mem[10922] = 126;
razn_h_mem[10923] = 2;
razn_h_mem[10924] = 132;
razn_h_mem[10925] = 8;
razn_h_mem[10926] = 138;
razn_h_mem[10927] = 14;
razn_h_mem[10928] = 144;
razn_h_mem[10929] = 20;
razn_h_mem[10930] = 150;
razn_h_mem[10931] = 26;
razn_h_mem[10932] = 156;
razn_h_mem[10933] = 32;
razn_h_mem[10934] = 162;
razn_h_mem[10935] = 38;
razn_h_mem[10936] = 168;
razn_h_mem[10937] = 44;
razn_h_mem[10938] = 174;
razn_h_mem[10939] = 50;
razn_h_mem[10940] = 180;
razn_h_mem[10941] = 56;
razn_h_mem[10942] = 186;
razn_h_mem[10943] = 62;
razn_h_mem[10944] = 192;
razn_h_mem[10945] = 68;
razn_h_mem[10946] = 198;
razn_h_mem[10947] = 74;
razn_h_mem[10948] = 204;
razn_h_mem[10949] = 80;
razn_h_mem[10950] = 210;
razn_h_mem[10951] = 86;
razn_h_mem[10952] = 216;
razn_h_mem[10953] = 92;
razn_h_mem[10954] = 222;
razn_h_mem[10955] = 98;
razn_h_mem[10956] = 228;
razn_h_mem[10957] = 104;
razn_h_mem[10958] = 234;
razn_h_mem[10959] = 110;
razn_h_mem[10960] = 240;
razn_h_mem[10961] = 116;
razn_h_mem[10962] = 246;
razn_h_mem[10963] = 122;
razn_h_mem[10964] = 252;
razn_h_mem[10965] = 128;
razn_h_mem[10966] = 4;
razn_h_mem[10967] = 134;
razn_h_mem[10968] = 10;
razn_h_mem[10969] = 140;
razn_h_mem[10970] = 16;
razn_h_mem[10971] = 146;
razn_h_mem[10972] = 22;
razn_h_mem[10973] = 152;
razn_h_mem[10974] = 28;
razn_h_mem[10975] = 158;
razn_h_mem[10976] = 34;
razn_h_mem[10977] = 164;
razn_h_mem[10978] = 40;
razn_h_mem[10979] = 170;
razn_h_mem[10980] = 46;
razn_h_mem[10981] = 176;
razn_h_mem[10982] = 52;
razn_h_mem[10983] = 182;
razn_h_mem[10984] = 58;
razn_h_mem[10985] = 188;
razn_h_mem[10986] = 64;
razn_h_mem[10987] = 194;
razn_h_mem[10988] = 70;
razn_h_mem[10989] = 200;
razn_h_mem[10990] = 76;
razn_h_mem[10991] = 206;
razn_h_mem[10992] = 82;
razn_h_mem[10993] = 212;
razn_h_mem[10994] = 88;
razn_h_mem[10995] = 218;
razn_h_mem[10996] = 94;
razn_h_mem[10997] = 224;
razn_h_mem[10998] = 100;
razn_h_mem[10999] = 230;
razn_h_mem[11000] = 106;
razn_h_mem[11001] = 236;
razn_h_mem[11002] = 112;
razn_h_mem[11003] = 242;
razn_h_mem[11004] = 118;
razn_h_mem[11005] = 248;
razn_h_mem[11006] = 124;
razn_h_mem[11007] = 255;
razn_h_mem[11008] = 0;
razn_h_mem[11009] = 130;
razn_h_mem[11010] = 6;
razn_h_mem[11011] = 136;
razn_h_mem[11012] = 12;
razn_h_mem[11013] = 142;
razn_h_mem[11014] = 18;
razn_h_mem[11015] = 148;
razn_h_mem[11016] = 24;
razn_h_mem[11017] = 154;
razn_h_mem[11018] = 30;
razn_h_mem[11019] = 160;
razn_h_mem[11020] = 36;
razn_h_mem[11021] = 166;
razn_h_mem[11022] = 42;
razn_h_mem[11023] = 172;
razn_h_mem[11024] = 48;
razn_h_mem[11025] = 178;
razn_h_mem[11026] = 54;
razn_h_mem[11027] = 184;
razn_h_mem[11028] = 60;
razn_h_mem[11029] = 190;
razn_h_mem[11030] = 66;
razn_h_mem[11031] = 196;
razn_h_mem[11032] = 72;
razn_h_mem[11033] = 202;
razn_h_mem[11034] = 78;
razn_h_mem[11035] = 208;
razn_h_mem[11036] = 84;
razn_h_mem[11037] = 214;
razn_h_mem[11038] = 90;
razn_h_mem[11039] = 220;
razn_h_mem[11040] = 96;
razn_h_mem[11041] = 226;
razn_h_mem[11042] = 102;
razn_h_mem[11043] = 232;
razn_h_mem[11044] = 108;
razn_h_mem[11045] = 238;
razn_h_mem[11046] = 114;
razn_h_mem[11047] = 244;
razn_h_mem[11048] = 120;
razn_h_mem[11049] = 250;
razn_h_mem[11050] = 126;
razn_h_mem[11051] = 2;
razn_h_mem[11052] = 132;
razn_h_mem[11053] = 8;
razn_h_mem[11054] = 138;
razn_h_mem[11055] = 14;
razn_h_mem[11056] = 144;
razn_h_mem[11057] = 20;
razn_h_mem[11058] = 150;
razn_h_mem[11059] = 26;
razn_h_mem[11060] = 156;
razn_h_mem[11061] = 32;
razn_h_mem[11062] = 162;
razn_h_mem[11063] = 38;
razn_h_mem[11064] = 168;
razn_h_mem[11065] = 44;
razn_h_mem[11066] = 174;
razn_h_mem[11067] = 50;
razn_h_mem[11068] = 180;
razn_h_mem[11069] = 56;
razn_h_mem[11070] = 186;
razn_h_mem[11071] = 62;
razn_h_mem[11072] = 192;
razn_h_mem[11073] = 68;
razn_h_mem[11074] = 198;
razn_h_mem[11075] = 74;
razn_h_mem[11076] = 204;
razn_h_mem[11077] = 80;
razn_h_mem[11078] = 210;
razn_h_mem[11079] = 86;
razn_h_mem[11080] = 216;
razn_h_mem[11081] = 92;
razn_h_mem[11082] = 222;
razn_h_mem[11083] = 98;
razn_h_mem[11084] = 228;
razn_h_mem[11085] = 104;
razn_h_mem[11086] = 234;
razn_h_mem[11087] = 110;
razn_h_mem[11088] = 240;
razn_h_mem[11089] = 116;
razn_h_mem[11090] = 246;
razn_h_mem[11091] = 122;
razn_h_mem[11092] = 252;
razn_h_mem[11093] = 128;
razn_h_mem[11094] = 4;
razn_h_mem[11095] = 134;
razn_h_mem[11096] = 10;
razn_h_mem[11097] = 140;
razn_h_mem[11098] = 16;
razn_h_mem[11099] = 146;
razn_h_mem[11100] = 22;
razn_h_mem[11101] = 152;
razn_h_mem[11102] = 28;
razn_h_mem[11103] = 158;
razn_h_mem[11104] = 34;
razn_h_mem[11105] = 164;
razn_h_mem[11106] = 40;
razn_h_mem[11107] = 170;
razn_h_mem[11108] = 46;
razn_h_mem[11109] = 176;
razn_h_mem[11110] = 52;
razn_h_mem[11111] = 182;
razn_h_mem[11112] = 58;
razn_h_mem[11113] = 188;
razn_h_mem[11114] = 64;
razn_h_mem[11115] = 194;
razn_h_mem[11116] = 70;
razn_h_mem[11117] = 200;
razn_h_mem[11118] = 76;
razn_h_mem[11119] = 206;
razn_h_mem[11120] = 82;
razn_h_mem[11121] = 212;
razn_h_mem[11122] = 88;
razn_h_mem[11123] = 218;
razn_h_mem[11124] = 94;
razn_h_mem[11125] = 224;
razn_h_mem[11126] = 100;
razn_h_mem[11127] = 230;
razn_h_mem[11128] = 106;
razn_h_mem[11129] = 236;
razn_h_mem[11130] = 112;
razn_h_mem[11131] = 242;
razn_h_mem[11132] = 118;
razn_h_mem[11133] = 248;
razn_h_mem[11134] = 124;
razn_h_mem[11135] = 255;
razn_h_mem[11136] = 0;
razn_h_mem[11137] = 130;
razn_h_mem[11138] = 6;
razn_h_mem[11139] = 136;
razn_h_mem[11140] = 12;
razn_h_mem[11141] = 142;
razn_h_mem[11142] = 18;
razn_h_mem[11143] = 148;
razn_h_mem[11144] = 24;
razn_h_mem[11145] = 154;
razn_h_mem[11146] = 30;
razn_h_mem[11147] = 160;
razn_h_mem[11148] = 36;
razn_h_mem[11149] = 166;
razn_h_mem[11150] = 42;
razn_h_mem[11151] = 172;
razn_h_mem[11152] = 48;
razn_h_mem[11153] = 178;
razn_h_mem[11154] = 54;
razn_h_mem[11155] = 184;
razn_h_mem[11156] = 60;
razn_h_mem[11157] = 190;
razn_h_mem[11158] = 66;
razn_h_mem[11159] = 196;
razn_h_mem[11160] = 72;
razn_h_mem[11161] = 202;
razn_h_mem[11162] = 78;
razn_h_mem[11163] = 208;
razn_h_mem[11164] = 84;
razn_h_mem[11165] = 214;
razn_h_mem[11166] = 90;
razn_h_mem[11167] = 220;
razn_h_mem[11168] = 96;
razn_h_mem[11169] = 226;
razn_h_mem[11170] = 102;
razn_h_mem[11171] = 232;
razn_h_mem[11172] = 108;
razn_h_mem[11173] = 238;
razn_h_mem[11174] = 114;
razn_h_mem[11175] = 244;
razn_h_mem[11176] = 120;
razn_h_mem[11177] = 250;
razn_h_mem[11178] = 126;
razn_h_mem[11179] = 2;
razn_h_mem[11180] = 132;
razn_h_mem[11181] = 8;
razn_h_mem[11182] = 138;
razn_h_mem[11183] = 14;
razn_h_mem[11184] = 144;
razn_h_mem[11185] = 20;
razn_h_mem[11186] = 150;
razn_h_mem[11187] = 26;
razn_h_mem[11188] = 156;
razn_h_mem[11189] = 32;
razn_h_mem[11190] = 162;
razn_h_mem[11191] = 38;
razn_h_mem[11192] = 168;
razn_h_mem[11193] = 44;
razn_h_mem[11194] = 174;
razn_h_mem[11195] = 50;
razn_h_mem[11196] = 180;
razn_h_mem[11197] = 56;
razn_h_mem[11198] = 186;
razn_h_mem[11199] = 62;
razn_h_mem[11200] = 192;
razn_h_mem[11201] = 68;
razn_h_mem[11202] = 198;
razn_h_mem[11203] = 74;
razn_h_mem[11204] = 204;
razn_h_mem[11205] = 80;
razn_h_mem[11206] = 210;
razn_h_mem[11207] = 86;
razn_h_mem[11208] = 216;
razn_h_mem[11209] = 92;
razn_h_mem[11210] = 222;
razn_h_mem[11211] = 98;
razn_h_mem[11212] = 228;
razn_h_mem[11213] = 104;
razn_h_mem[11214] = 234;
razn_h_mem[11215] = 110;
razn_h_mem[11216] = 240;
razn_h_mem[11217] = 116;
razn_h_mem[11218] = 246;
razn_h_mem[11219] = 122;
razn_h_mem[11220] = 252;
razn_h_mem[11221] = 128;
razn_h_mem[11222] = 4;
razn_h_mem[11223] = 134;
razn_h_mem[11224] = 10;
razn_h_mem[11225] = 140;
razn_h_mem[11226] = 16;
razn_h_mem[11227] = 146;
razn_h_mem[11228] = 22;
razn_h_mem[11229] = 152;
razn_h_mem[11230] = 28;
razn_h_mem[11231] = 158;
razn_h_mem[11232] = 34;
razn_h_mem[11233] = 164;
razn_h_mem[11234] = 40;
razn_h_mem[11235] = 170;
razn_h_mem[11236] = 46;
razn_h_mem[11237] = 176;
razn_h_mem[11238] = 52;
razn_h_mem[11239] = 182;
razn_h_mem[11240] = 58;
razn_h_mem[11241] = 188;
razn_h_mem[11242] = 64;
razn_h_mem[11243] = 194;
razn_h_mem[11244] = 70;
razn_h_mem[11245] = 200;
razn_h_mem[11246] = 76;
razn_h_mem[11247] = 206;
razn_h_mem[11248] = 82;
razn_h_mem[11249] = 212;
razn_h_mem[11250] = 88;
razn_h_mem[11251] = 218;
razn_h_mem[11252] = 94;
razn_h_mem[11253] = 224;
razn_h_mem[11254] = 100;
razn_h_mem[11255] = 230;
razn_h_mem[11256] = 106;
razn_h_mem[11257] = 236;
razn_h_mem[11258] = 112;
razn_h_mem[11259] = 242;
razn_h_mem[11260] = 118;
razn_h_mem[11261] = 248;
razn_h_mem[11262] = 124;
razn_h_mem[11263] = 255;
razn_h_mem[11264] = 0;
razn_h_mem[11265] = 130;
razn_h_mem[11266] = 6;
razn_h_mem[11267] = 136;
razn_h_mem[11268] = 12;
razn_h_mem[11269] = 142;
razn_h_mem[11270] = 18;
razn_h_mem[11271] = 148;
razn_h_mem[11272] = 24;
razn_h_mem[11273] = 154;
razn_h_mem[11274] = 30;
razn_h_mem[11275] = 160;
razn_h_mem[11276] = 36;
razn_h_mem[11277] = 166;
razn_h_mem[11278] = 42;
razn_h_mem[11279] = 172;
razn_h_mem[11280] = 48;
razn_h_mem[11281] = 178;
razn_h_mem[11282] = 54;
razn_h_mem[11283] = 184;
razn_h_mem[11284] = 60;
razn_h_mem[11285] = 190;
razn_h_mem[11286] = 66;
razn_h_mem[11287] = 196;
razn_h_mem[11288] = 72;
razn_h_mem[11289] = 202;
razn_h_mem[11290] = 78;
razn_h_mem[11291] = 208;
razn_h_mem[11292] = 84;
razn_h_mem[11293] = 214;
razn_h_mem[11294] = 90;
razn_h_mem[11295] = 220;
razn_h_mem[11296] = 96;
razn_h_mem[11297] = 226;
razn_h_mem[11298] = 102;
razn_h_mem[11299] = 232;
razn_h_mem[11300] = 108;
razn_h_mem[11301] = 238;
razn_h_mem[11302] = 114;
razn_h_mem[11303] = 244;
razn_h_mem[11304] = 120;
razn_h_mem[11305] = 250;
razn_h_mem[11306] = 126;
razn_h_mem[11307] = 2;
razn_h_mem[11308] = 132;
razn_h_mem[11309] = 8;
razn_h_mem[11310] = 138;
razn_h_mem[11311] = 14;
razn_h_mem[11312] = 144;
razn_h_mem[11313] = 20;
razn_h_mem[11314] = 150;
razn_h_mem[11315] = 26;
razn_h_mem[11316] = 156;
razn_h_mem[11317] = 32;
razn_h_mem[11318] = 162;
razn_h_mem[11319] = 38;
razn_h_mem[11320] = 168;
razn_h_mem[11321] = 44;
razn_h_mem[11322] = 174;
razn_h_mem[11323] = 50;
razn_h_mem[11324] = 180;
razn_h_mem[11325] = 56;
razn_h_mem[11326] = 186;
razn_h_mem[11327] = 62;
razn_h_mem[11328] = 192;
razn_h_mem[11329] = 68;
razn_h_mem[11330] = 198;
razn_h_mem[11331] = 74;
razn_h_mem[11332] = 204;
razn_h_mem[11333] = 80;
razn_h_mem[11334] = 210;
razn_h_mem[11335] = 86;
razn_h_mem[11336] = 216;
razn_h_mem[11337] = 92;
razn_h_mem[11338] = 222;
razn_h_mem[11339] = 98;
razn_h_mem[11340] = 228;
razn_h_mem[11341] = 104;
razn_h_mem[11342] = 234;
razn_h_mem[11343] = 110;
razn_h_mem[11344] = 240;
razn_h_mem[11345] = 116;
razn_h_mem[11346] = 246;
razn_h_mem[11347] = 122;
razn_h_mem[11348] = 252;
razn_h_mem[11349] = 128;
razn_h_mem[11350] = 4;
razn_h_mem[11351] = 134;
razn_h_mem[11352] = 10;
razn_h_mem[11353] = 140;
razn_h_mem[11354] = 16;
razn_h_mem[11355] = 146;
razn_h_mem[11356] = 22;
razn_h_mem[11357] = 152;
razn_h_mem[11358] = 28;
razn_h_mem[11359] = 158;
razn_h_mem[11360] = 34;
razn_h_mem[11361] = 164;
razn_h_mem[11362] = 40;
razn_h_mem[11363] = 170;
razn_h_mem[11364] = 46;
razn_h_mem[11365] = 176;
razn_h_mem[11366] = 52;
razn_h_mem[11367] = 182;
razn_h_mem[11368] = 58;
razn_h_mem[11369] = 188;
razn_h_mem[11370] = 64;
razn_h_mem[11371] = 194;
razn_h_mem[11372] = 70;
razn_h_mem[11373] = 200;
razn_h_mem[11374] = 76;
razn_h_mem[11375] = 206;
razn_h_mem[11376] = 82;
razn_h_mem[11377] = 212;
razn_h_mem[11378] = 88;
razn_h_mem[11379] = 218;
razn_h_mem[11380] = 94;
razn_h_mem[11381] = 224;
razn_h_mem[11382] = 100;
razn_h_mem[11383] = 230;
razn_h_mem[11384] = 106;
razn_h_mem[11385] = 236;
razn_h_mem[11386] = 112;
razn_h_mem[11387] = 242;
razn_h_mem[11388] = 118;
razn_h_mem[11389] = 248;
razn_h_mem[11390] = 124;
razn_h_mem[11391] = 255;
razn_h_mem[11392] = 0;
razn_h_mem[11393] = 130;
razn_h_mem[11394] = 6;
razn_h_mem[11395] = 136;
razn_h_mem[11396] = 12;
razn_h_mem[11397] = 142;
razn_h_mem[11398] = 18;
razn_h_mem[11399] = 148;
razn_h_mem[11400] = 24;
razn_h_mem[11401] = 154;
razn_h_mem[11402] = 30;
razn_h_mem[11403] = 160;
razn_h_mem[11404] = 36;
razn_h_mem[11405] = 166;
razn_h_mem[11406] = 42;
razn_h_mem[11407] = 172;
razn_h_mem[11408] = 48;
razn_h_mem[11409] = 178;
razn_h_mem[11410] = 54;
razn_h_mem[11411] = 184;
razn_h_mem[11412] = 60;
razn_h_mem[11413] = 190;
razn_h_mem[11414] = 66;
razn_h_mem[11415] = 196;
razn_h_mem[11416] = 72;
razn_h_mem[11417] = 202;
razn_h_mem[11418] = 78;
razn_h_mem[11419] = 208;
razn_h_mem[11420] = 84;
razn_h_mem[11421] = 214;
razn_h_mem[11422] = 90;
razn_h_mem[11423] = 220;
razn_h_mem[11424] = 96;
razn_h_mem[11425] = 226;
razn_h_mem[11426] = 102;
razn_h_mem[11427] = 232;
razn_h_mem[11428] = 108;
razn_h_mem[11429] = 238;
razn_h_mem[11430] = 114;
razn_h_mem[11431] = 244;
razn_h_mem[11432] = 120;
razn_h_mem[11433] = 250;
razn_h_mem[11434] = 126;
razn_h_mem[11435] = 2;
razn_h_mem[11436] = 132;
razn_h_mem[11437] = 8;
razn_h_mem[11438] = 138;
razn_h_mem[11439] = 14;
razn_h_mem[11440] = 144;
razn_h_mem[11441] = 20;
razn_h_mem[11442] = 150;
razn_h_mem[11443] = 26;
razn_h_mem[11444] = 156;
razn_h_mem[11445] = 32;
razn_h_mem[11446] = 162;
razn_h_mem[11447] = 38;
razn_h_mem[11448] = 168;
razn_h_mem[11449] = 44;
razn_h_mem[11450] = 174;
razn_h_mem[11451] = 50;
razn_h_mem[11452] = 180;
razn_h_mem[11453] = 56;
razn_h_mem[11454] = 186;
razn_h_mem[11455] = 62;
razn_h_mem[11456] = 192;
razn_h_mem[11457] = 68;
razn_h_mem[11458] = 198;
razn_h_mem[11459] = 74;
razn_h_mem[11460] = 204;
razn_h_mem[11461] = 80;
razn_h_mem[11462] = 210;
razn_h_mem[11463] = 86;
razn_h_mem[11464] = 216;
razn_h_mem[11465] = 92;
razn_h_mem[11466] = 222;
razn_h_mem[11467] = 98;
razn_h_mem[11468] = 228;
razn_h_mem[11469] = 104;
razn_h_mem[11470] = 234;
razn_h_mem[11471] = 110;
razn_h_mem[11472] = 240;
razn_h_mem[11473] = 116;
razn_h_mem[11474] = 246;
razn_h_mem[11475] = 122;
razn_h_mem[11476] = 252;
razn_h_mem[11477] = 128;
razn_h_mem[11478] = 4;
razn_h_mem[11479] = 134;
razn_h_mem[11480] = 10;
razn_h_mem[11481] = 140;
razn_h_mem[11482] = 16;
razn_h_mem[11483] = 146;
razn_h_mem[11484] = 22;
razn_h_mem[11485] = 152;
razn_h_mem[11486] = 28;
razn_h_mem[11487] = 158;
razn_h_mem[11488] = 34;
razn_h_mem[11489] = 164;
razn_h_mem[11490] = 40;
razn_h_mem[11491] = 170;
razn_h_mem[11492] = 46;
razn_h_mem[11493] = 176;
razn_h_mem[11494] = 52;
razn_h_mem[11495] = 182;
razn_h_mem[11496] = 58;
razn_h_mem[11497] = 188;
razn_h_mem[11498] = 64;
razn_h_mem[11499] = 194;
razn_h_mem[11500] = 70;
razn_h_mem[11501] = 200;
razn_h_mem[11502] = 76;
razn_h_mem[11503] = 206;
razn_h_mem[11504] = 82;
razn_h_mem[11505] = 212;
razn_h_mem[11506] = 88;
razn_h_mem[11507] = 218;
razn_h_mem[11508] = 94;
razn_h_mem[11509] = 224;
razn_h_mem[11510] = 100;
razn_h_mem[11511] = 230;
razn_h_mem[11512] = 106;
razn_h_mem[11513] = 236;
razn_h_mem[11514] = 112;
razn_h_mem[11515] = 242;
razn_h_mem[11516] = 118;
razn_h_mem[11517] = 248;
razn_h_mem[11518] = 124;
razn_h_mem[11519] = 255;
razn_h_mem[11520] = 0;
razn_h_mem[11521] = 130;
razn_h_mem[11522] = 6;
razn_h_mem[11523] = 136;
razn_h_mem[11524] = 12;
razn_h_mem[11525] = 142;
razn_h_mem[11526] = 18;
razn_h_mem[11527] = 148;
razn_h_mem[11528] = 24;
razn_h_mem[11529] = 154;
razn_h_mem[11530] = 30;
razn_h_mem[11531] = 160;
razn_h_mem[11532] = 36;
razn_h_mem[11533] = 166;
razn_h_mem[11534] = 42;
razn_h_mem[11535] = 172;
razn_h_mem[11536] = 48;
razn_h_mem[11537] = 178;
razn_h_mem[11538] = 54;
razn_h_mem[11539] = 184;
razn_h_mem[11540] = 60;
razn_h_mem[11541] = 190;
razn_h_mem[11542] = 66;
razn_h_mem[11543] = 196;
razn_h_mem[11544] = 72;
razn_h_mem[11545] = 202;
razn_h_mem[11546] = 78;
razn_h_mem[11547] = 208;
razn_h_mem[11548] = 84;
razn_h_mem[11549] = 214;
razn_h_mem[11550] = 90;
razn_h_mem[11551] = 220;
razn_h_mem[11552] = 96;
razn_h_mem[11553] = 226;
razn_h_mem[11554] = 102;
razn_h_mem[11555] = 232;
razn_h_mem[11556] = 108;
razn_h_mem[11557] = 238;
razn_h_mem[11558] = 114;
razn_h_mem[11559] = 244;
razn_h_mem[11560] = 120;
razn_h_mem[11561] = 250;
razn_h_mem[11562] = 126;
razn_h_mem[11563] = 2;
razn_h_mem[11564] = 132;
razn_h_mem[11565] = 8;
razn_h_mem[11566] = 138;
razn_h_mem[11567] = 14;
razn_h_mem[11568] = 144;
razn_h_mem[11569] = 20;
razn_h_mem[11570] = 150;
razn_h_mem[11571] = 26;
razn_h_mem[11572] = 156;
razn_h_mem[11573] = 32;
razn_h_mem[11574] = 162;
razn_h_mem[11575] = 38;
razn_h_mem[11576] = 168;
razn_h_mem[11577] = 44;
razn_h_mem[11578] = 174;
razn_h_mem[11579] = 50;
razn_h_mem[11580] = 180;
razn_h_mem[11581] = 56;
razn_h_mem[11582] = 186;
razn_h_mem[11583] = 62;
razn_h_mem[11584] = 192;
razn_h_mem[11585] = 68;
razn_h_mem[11586] = 198;
razn_h_mem[11587] = 74;
razn_h_mem[11588] = 204;
razn_h_mem[11589] = 80;
razn_h_mem[11590] = 210;
razn_h_mem[11591] = 86;
razn_h_mem[11592] = 216;
razn_h_mem[11593] = 92;
razn_h_mem[11594] = 222;
razn_h_mem[11595] = 98;
razn_h_mem[11596] = 228;
razn_h_mem[11597] = 104;
razn_h_mem[11598] = 234;
razn_h_mem[11599] = 110;
razn_h_mem[11600] = 240;
razn_h_mem[11601] = 116;
razn_h_mem[11602] = 246;
razn_h_mem[11603] = 122;
razn_h_mem[11604] = 252;
razn_h_mem[11605] = 128;
razn_h_mem[11606] = 4;
razn_h_mem[11607] = 134;
razn_h_mem[11608] = 10;
razn_h_mem[11609] = 140;
razn_h_mem[11610] = 16;
razn_h_mem[11611] = 146;
razn_h_mem[11612] = 22;
razn_h_mem[11613] = 152;
razn_h_mem[11614] = 28;
razn_h_mem[11615] = 158;
razn_h_mem[11616] = 34;
razn_h_mem[11617] = 164;
razn_h_mem[11618] = 40;
razn_h_mem[11619] = 170;
razn_h_mem[11620] = 46;
razn_h_mem[11621] = 176;
razn_h_mem[11622] = 52;
razn_h_mem[11623] = 182;
razn_h_mem[11624] = 58;
razn_h_mem[11625] = 188;
razn_h_mem[11626] = 64;
razn_h_mem[11627] = 194;
razn_h_mem[11628] = 70;
razn_h_mem[11629] = 200;
razn_h_mem[11630] = 76;
razn_h_mem[11631] = 206;
razn_h_mem[11632] = 82;
razn_h_mem[11633] = 212;
razn_h_mem[11634] = 88;
razn_h_mem[11635] = 218;
razn_h_mem[11636] = 94;
razn_h_mem[11637] = 224;
razn_h_mem[11638] = 100;
razn_h_mem[11639] = 230;
razn_h_mem[11640] = 106;
razn_h_mem[11641] = 236;
razn_h_mem[11642] = 112;
razn_h_mem[11643] = 242;
razn_h_mem[11644] = 118;
razn_h_mem[11645] = 248;
razn_h_mem[11646] = 124;
razn_h_mem[11647] = 255;
razn_h_mem[11648] = 0;
razn_h_mem[11649] = 130;
razn_h_mem[11650] = 6;
razn_h_mem[11651] = 136;
razn_h_mem[11652] = 12;
razn_h_mem[11653] = 142;
razn_h_mem[11654] = 18;
razn_h_mem[11655] = 148;
razn_h_mem[11656] = 24;
razn_h_mem[11657] = 154;
razn_h_mem[11658] = 30;
razn_h_mem[11659] = 160;
razn_h_mem[11660] = 36;
razn_h_mem[11661] = 166;
razn_h_mem[11662] = 42;
razn_h_mem[11663] = 172;
razn_h_mem[11664] = 48;
razn_h_mem[11665] = 178;
razn_h_mem[11666] = 54;
razn_h_mem[11667] = 184;
razn_h_mem[11668] = 60;
razn_h_mem[11669] = 190;
razn_h_mem[11670] = 66;
razn_h_mem[11671] = 196;
razn_h_mem[11672] = 72;
razn_h_mem[11673] = 202;
razn_h_mem[11674] = 78;
razn_h_mem[11675] = 208;
razn_h_mem[11676] = 84;
razn_h_mem[11677] = 214;
razn_h_mem[11678] = 90;
razn_h_mem[11679] = 220;
razn_h_mem[11680] = 96;
razn_h_mem[11681] = 226;
razn_h_mem[11682] = 102;
razn_h_mem[11683] = 232;
razn_h_mem[11684] = 108;
razn_h_mem[11685] = 238;
razn_h_mem[11686] = 114;
razn_h_mem[11687] = 244;
razn_h_mem[11688] = 120;
razn_h_mem[11689] = 250;
razn_h_mem[11690] = 126;
razn_h_mem[11691] = 2;
razn_h_mem[11692] = 132;
razn_h_mem[11693] = 8;
razn_h_mem[11694] = 138;
razn_h_mem[11695] = 14;
razn_h_mem[11696] = 144;
razn_h_mem[11697] = 20;
razn_h_mem[11698] = 150;
razn_h_mem[11699] = 26;
razn_h_mem[11700] = 156;
razn_h_mem[11701] = 32;
razn_h_mem[11702] = 162;
razn_h_mem[11703] = 38;
razn_h_mem[11704] = 168;
razn_h_mem[11705] = 44;
razn_h_mem[11706] = 174;
razn_h_mem[11707] = 50;
razn_h_mem[11708] = 180;
razn_h_mem[11709] = 56;
razn_h_mem[11710] = 186;
razn_h_mem[11711] = 62;
razn_h_mem[11712] = 192;
razn_h_mem[11713] = 68;
razn_h_mem[11714] = 198;
razn_h_mem[11715] = 74;
razn_h_mem[11716] = 204;
razn_h_mem[11717] = 80;
razn_h_mem[11718] = 210;
razn_h_mem[11719] = 86;
razn_h_mem[11720] = 216;
razn_h_mem[11721] = 92;
razn_h_mem[11722] = 222;
razn_h_mem[11723] = 98;
razn_h_mem[11724] = 228;
razn_h_mem[11725] = 104;
razn_h_mem[11726] = 234;
razn_h_mem[11727] = 110;
razn_h_mem[11728] = 240;
razn_h_mem[11729] = 116;
razn_h_mem[11730] = 246;
razn_h_mem[11731] = 122;
razn_h_mem[11732] = 252;
razn_h_mem[11733] = 128;
razn_h_mem[11734] = 4;
razn_h_mem[11735] = 134;
razn_h_mem[11736] = 10;
razn_h_mem[11737] = 140;
razn_h_mem[11738] = 16;
razn_h_mem[11739] = 146;
razn_h_mem[11740] = 22;
razn_h_mem[11741] = 152;
razn_h_mem[11742] = 28;
razn_h_mem[11743] = 158;
razn_h_mem[11744] = 34;
razn_h_mem[11745] = 164;
razn_h_mem[11746] = 40;
razn_h_mem[11747] = 170;
razn_h_mem[11748] = 46;
razn_h_mem[11749] = 176;
razn_h_mem[11750] = 52;
razn_h_mem[11751] = 182;
razn_h_mem[11752] = 58;
razn_h_mem[11753] = 188;
razn_h_mem[11754] = 64;
razn_h_mem[11755] = 194;
razn_h_mem[11756] = 70;
razn_h_mem[11757] = 200;
razn_h_mem[11758] = 76;
razn_h_mem[11759] = 206;
razn_h_mem[11760] = 82;
razn_h_mem[11761] = 212;
razn_h_mem[11762] = 88;
razn_h_mem[11763] = 218;
razn_h_mem[11764] = 94;
razn_h_mem[11765] = 224;
razn_h_mem[11766] = 100;
razn_h_mem[11767] = 230;
razn_h_mem[11768] = 106;
razn_h_mem[11769] = 236;
razn_h_mem[11770] = 112;
razn_h_mem[11771] = 242;
razn_h_mem[11772] = 118;
razn_h_mem[11773] = 248;
razn_h_mem[11774] = 124;
razn_h_mem[11775] = 255;
razn_h_mem[11776] = 0;
razn_h_mem[11777] = 130;
razn_h_mem[11778] = 6;
razn_h_mem[11779] = 136;
razn_h_mem[11780] = 12;
razn_h_mem[11781] = 142;
razn_h_mem[11782] = 18;
razn_h_mem[11783] = 148;
razn_h_mem[11784] = 24;
razn_h_mem[11785] = 154;
razn_h_mem[11786] = 30;
razn_h_mem[11787] = 160;
razn_h_mem[11788] = 36;
razn_h_mem[11789] = 166;
razn_h_mem[11790] = 42;
razn_h_mem[11791] = 172;
razn_h_mem[11792] = 48;
razn_h_mem[11793] = 178;
razn_h_mem[11794] = 54;
razn_h_mem[11795] = 184;
razn_h_mem[11796] = 60;
razn_h_mem[11797] = 190;
razn_h_mem[11798] = 66;
razn_h_mem[11799] = 196;
razn_h_mem[11800] = 72;
razn_h_mem[11801] = 202;
razn_h_mem[11802] = 78;
razn_h_mem[11803] = 208;
razn_h_mem[11804] = 84;
razn_h_mem[11805] = 214;
razn_h_mem[11806] = 90;
razn_h_mem[11807] = 220;
razn_h_mem[11808] = 96;
razn_h_mem[11809] = 226;
razn_h_mem[11810] = 102;
razn_h_mem[11811] = 232;
razn_h_mem[11812] = 108;
razn_h_mem[11813] = 238;
razn_h_mem[11814] = 114;
razn_h_mem[11815] = 244;
razn_h_mem[11816] = 120;
razn_h_mem[11817] = 250;
razn_h_mem[11818] = 126;
razn_h_mem[11819] = 2;
razn_h_mem[11820] = 132;
razn_h_mem[11821] = 8;
razn_h_mem[11822] = 138;
razn_h_mem[11823] = 14;
razn_h_mem[11824] = 144;
razn_h_mem[11825] = 20;
razn_h_mem[11826] = 150;
razn_h_mem[11827] = 26;
razn_h_mem[11828] = 156;
razn_h_mem[11829] = 32;
razn_h_mem[11830] = 162;
razn_h_mem[11831] = 38;
razn_h_mem[11832] = 168;
razn_h_mem[11833] = 44;
razn_h_mem[11834] = 174;
razn_h_mem[11835] = 50;
razn_h_mem[11836] = 180;
razn_h_mem[11837] = 56;
razn_h_mem[11838] = 186;
razn_h_mem[11839] = 62;
razn_h_mem[11840] = 192;
razn_h_mem[11841] = 68;
razn_h_mem[11842] = 198;
razn_h_mem[11843] = 74;
razn_h_mem[11844] = 204;
razn_h_mem[11845] = 80;
razn_h_mem[11846] = 210;
razn_h_mem[11847] = 86;
razn_h_mem[11848] = 216;
razn_h_mem[11849] = 92;
razn_h_mem[11850] = 222;
razn_h_mem[11851] = 98;
razn_h_mem[11852] = 228;
razn_h_mem[11853] = 104;
razn_h_mem[11854] = 234;
razn_h_mem[11855] = 110;
razn_h_mem[11856] = 240;
razn_h_mem[11857] = 116;
razn_h_mem[11858] = 246;
razn_h_mem[11859] = 122;
razn_h_mem[11860] = 252;
razn_h_mem[11861] = 128;
razn_h_mem[11862] = 4;
razn_h_mem[11863] = 134;
razn_h_mem[11864] = 10;
razn_h_mem[11865] = 140;
razn_h_mem[11866] = 16;
razn_h_mem[11867] = 146;
razn_h_mem[11868] = 22;
razn_h_mem[11869] = 152;
razn_h_mem[11870] = 28;
razn_h_mem[11871] = 158;
razn_h_mem[11872] = 34;
razn_h_mem[11873] = 164;
razn_h_mem[11874] = 40;
razn_h_mem[11875] = 170;
razn_h_mem[11876] = 46;
razn_h_mem[11877] = 176;
razn_h_mem[11878] = 52;
razn_h_mem[11879] = 182;
razn_h_mem[11880] = 58;
razn_h_mem[11881] = 188;
razn_h_mem[11882] = 64;
razn_h_mem[11883] = 194;
razn_h_mem[11884] = 70;
razn_h_mem[11885] = 200;
razn_h_mem[11886] = 76;
razn_h_mem[11887] = 206;
razn_h_mem[11888] = 82;
razn_h_mem[11889] = 212;
razn_h_mem[11890] = 88;
razn_h_mem[11891] = 218;
razn_h_mem[11892] = 94;
razn_h_mem[11893] = 224;
razn_h_mem[11894] = 100;
razn_h_mem[11895] = 230;
razn_h_mem[11896] = 106;
razn_h_mem[11897] = 236;
razn_h_mem[11898] = 112;
razn_h_mem[11899] = 242;
razn_h_mem[11900] = 118;
razn_h_mem[11901] = 248;
razn_h_mem[11902] = 124;
razn_h_mem[11903] = 255;
razn_h_mem[11904] = 0;
razn_h_mem[11905] = 130;
razn_h_mem[11906] = 6;
razn_h_mem[11907] = 136;
razn_h_mem[11908] = 12;
razn_h_mem[11909] = 142;
razn_h_mem[11910] = 18;
razn_h_mem[11911] = 148;
razn_h_mem[11912] = 24;
razn_h_mem[11913] = 154;
razn_h_mem[11914] = 30;
razn_h_mem[11915] = 160;
razn_h_mem[11916] = 36;
razn_h_mem[11917] = 166;
razn_h_mem[11918] = 42;
razn_h_mem[11919] = 172;
razn_h_mem[11920] = 48;
razn_h_mem[11921] = 178;
razn_h_mem[11922] = 54;
razn_h_mem[11923] = 184;
razn_h_mem[11924] = 60;
razn_h_mem[11925] = 190;
razn_h_mem[11926] = 66;
razn_h_mem[11927] = 196;
razn_h_mem[11928] = 72;
razn_h_mem[11929] = 202;
razn_h_mem[11930] = 78;
razn_h_mem[11931] = 208;
razn_h_mem[11932] = 84;
razn_h_mem[11933] = 214;
razn_h_mem[11934] = 90;
razn_h_mem[11935] = 220;
razn_h_mem[11936] = 96;
razn_h_mem[11937] = 226;
razn_h_mem[11938] = 102;
razn_h_mem[11939] = 232;
razn_h_mem[11940] = 108;
razn_h_mem[11941] = 238;
razn_h_mem[11942] = 114;
razn_h_mem[11943] = 244;
razn_h_mem[11944] = 120;
razn_h_mem[11945] = 250;
razn_h_mem[11946] = 126;
razn_h_mem[11947] = 2;
razn_h_mem[11948] = 132;
razn_h_mem[11949] = 8;
razn_h_mem[11950] = 138;
razn_h_mem[11951] = 14;
razn_h_mem[11952] = 144;
razn_h_mem[11953] = 20;
razn_h_mem[11954] = 150;
razn_h_mem[11955] = 26;
razn_h_mem[11956] = 156;
razn_h_mem[11957] = 32;
razn_h_mem[11958] = 162;
razn_h_mem[11959] = 38;
razn_h_mem[11960] = 168;
razn_h_mem[11961] = 44;
razn_h_mem[11962] = 174;
razn_h_mem[11963] = 50;
razn_h_mem[11964] = 180;
razn_h_mem[11965] = 56;
razn_h_mem[11966] = 186;
razn_h_mem[11967] = 62;
razn_h_mem[11968] = 192;
razn_h_mem[11969] = 68;
razn_h_mem[11970] = 198;
razn_h_mem[11971] = 74;
razn_h_mem[11972] = 204;
razn_h_mem[11973] = 80;
razn_h_mem[11974] = 210;
razn_h_mem[11975] = 86;
razn_h_mem[11976] = 216;
razn_h_mem[11977] = 92;
razn_h_mem[11978] = 222;
razn_h_mem[11979] = 98;
razn_h_mem[11980] = 228;
razn_h_mem[11981] = 104;
razn_h_mem[11982] = 234;
razn_h_mem[11983] = 110;
razn_h_mem[11984] = 240;
razn_h_mem[11985] = 116;
razn_h_mem[11986] = 246;
razn_h_mem[11987] = 122;
razn_h_mem[11988] = 252;
razn_h_mem[11989] = 128;
razn_h_mem[11990] = 4;
razn_h_mem[11991] = 134;
razn_h_mem[11992] = 10;
razn_h_mem[11993] = 140;
razn_h_mem[11994] = 16;
razn_h_mem[11995] = 146;
razn_h_mem[11996] = 22;
razn_h_mem[11997] = 152;
razn_h_mem[11998] = 28;
razn_h_mem[11999] = 158;
razn_h_mem[12000] = 34;
razn_h_mem[12001] = 164;
razn_h_mem[12002] = 40;
razn_h_mem[12003] = 170;
razn_h_mem[12004] = 46;
razn_h_mem[12005] = 176;
razn_h_mem[12006] = 52;
razn_h_mem[12007] = 182;
razn_h_mem[12008] = 58;
razn_h_mem[12009] = 188;
razn_h_mem[12010] = 64;
razn_h_mem[12011] = 194;
razn_h_mem[12012] = 70;
razn_h_mem[12013] = 200;
razn_h_mem[12014] = 76;
razn_h_mem[12015] = 206;
razn_h_mem[12016] = 82;
razn_h_mem[12017] = 212;
razn_h_mem[12018] = 88;
razn_h_mem[12019] = 218;
razn_h_mem[12020] = 94;
razn_h_mem[12021] = 224;
razn_h_mem[12022] = 100;
razn_h_mem[12023] = 230;
razn_h_mem[12024] = 106;
razn_h_mem[12025] = 236;
razn_h_mem[12026] = 112;
razn_h_mem[12027] = 242;
razn_h_mem[12028] = 118;
razn_h_mem[12029] = 248;
razn_h_mem[12030] = 124;
razn_h_mem[12031] = 255;
razn_h_mem[12032] = 0;
razn_h_mem[12033] = 130;
razn_h_mem[12034] = 6;
razn_h_mem[12035] = 136;
razn_h_mem[12036] = 12;
razn_h_mem[12037] = 142;
razn_h_mem[12038] = 18;
razn_h_mem[12039] = 148;
razn_h_mem[12040] = 24;
razn_h_mem[12041] = 154;
razn_h_mem[12042] = 30;
razn_h_mem[12043] = 160;
razn_h_mem[12044] = 36;
razn_h_mem[12045] = 166;
razn_h_mem[12046] = 42;
razn_h_mem[12047] = 172;
razn_h_mem[12048] = 48;
razn_h_mem[12049] = 178;
razn_h_mem[12050] = 54;
razn_h_mem[12051] = 184;
razn_h_mem[12052] = 60;
razn_h_mem[12053] = 190;
razn_h_mem[12054] = 66;
razn_h_mem[12055] = 196;
razn_h_mem[12056] = 72;
razn_h_mem[12057] = 202;
razn_h_mem[12058] = 78;
razn_h_mem[12059] = 208;
razn_h_mem[12060] = 84;
razn_h_mem[12061] = 214;
razn_h_mem[12062] = 90;
razn_h_mem[12063] = 220;
razn_h_mem[12064] = 96;
razn_h_mem[12065] = 226;
razn_h_mem[12066] = 102;
razn_h_mem[12067] = 232;
razn_h_mem[12068] = 108;
razn_h_mem[12069] = 238;
razn_h_mem[12070] = 114;
razn_h_mem[12071] = 244;
razn_h_mem[12072] = 120;
razn_h_mem[12073] = 250;
razn_h_mem[12074] = 126;
razn_h_mem[12075] = 2;
razn_h_mem[12076] = 132;
razn_h_mem[12077] = 8;
razn_h_mem[12078] = 138;
razn_h_mem[12079] = 14;
razn_h_mem[12080] = 144;
razn_h_mem[12081] = 20;
razn_h_mem[12082] = 150;
razn_h_mem[12083] = 26;
razn_h_mem[12084] = 156;
razn_h_mem[12085] = 32;
razn_h_mem[12086] = 162;
razn_h_mem[12087] = 38;
razn_h_mem[12088] = 168;
razn_h_mem[12089] = 44;
razn_h_mem[12090] = 174;
razn_h_mem[12091] = 50;
razn_h_mem[12092] = 180;
razn_h_mem[12093] = 56;
razn_h_mem[12094] = 186;
razn_h_mem[12095] = 62;
razn_h_mem[12096] = 192;
razn_h_mem[12097] = 68;
razn_h_mem[12098] = 198;
razn_h_mem[12099] = 74;
razn_h_mem[12100] = 204;
razn_h_mem[12101] = 80;
razn_h_mem[12102] = 210;
razn_h_mem[12103] = 86;
razn_h_mem[12104] = 216;
razn_h_mem[12105] = 92;
razn_h_mem[12106] = 222;
razn_h_mem[12107] = 98;
razn_h_mem[12108] = 228;
razn_h_mem[12109] = 104;
razn_h_mem[12110] = 234;
razn_h_mem[12111] = 110;
razn_h_mem[12112] = 240;
razn_h_mem[12113] = 116;
razn_h_mem[12114] = 246;
razn_h_mem[12115] = 122;
razn_h_mem[12116] = 252;
razn_h_mem[12117] = 128;
razn_h_mem[12118] = 4;
razn_h_mem[12119] = 134;
razn_h_mem[12120] = 10;
razn_h_mem[12121] = 140;
razn_h_mem[12122] = 16;
razn_h_mem[12123] = 146;
razn_h_mem[12124] = 22;
razn_h_mem[12125] = 152;
razn_h_mem[12126] = 28;
razn_h_mem[12127] = 158;
razn_h_mem[12128] = 34;
razn_h_mem[12129] = 164;
razn_h_mem[12130] = 40;
razn_h_mem[12131] = 170;
razn_h_mem[12132] = 46;
razn_h_mem[12133] = 176;
razn_h_mem[12134] = 52;
razn_h_mem[12135] = 182;
razn_h_mem[12136] = 58;
razn_h_mem[12137] = 188;
razn_h_mem[12138] = 64;
razn_h_mem[12139] = 194;
razn_h_mem[12140] = 70;
razn_h_mem[12141] = 200;
razn_h_mem[12142] = 76;
razn_h_mem[12143] = 206;
razn_h_mem[12144] = 82;
razn_h_mem[12145] = 212;
razn_h_mem[12146] = 88;
razn_h_mem[12147] = 218;
razn_h_mem[12148] = 94;
razn_h_mem[12149] = 224;
razn_h_mem[12150] = 100;
razn_h_mem[12151] = 230;
razn_h_mem[12152] = 106;
razn_h_mem[12153] = 236;
razn_h_mem[12154] = 112;
razn_h_mem[12155] = 242;
razn_h_mem[12156] = 118;
razn_h_mem[12157] = 248;
razn_h_mem[12158] = 124;
razn_h_mem[12159] = 255;
razn_h_mem[12160] = 0;
razn_h_mem[12161] = 130;
razn_h_mem[12162] = 6;
razn_h_mem[12163] = 136;
razn_h_mem[12164] = 12;
razn_h_mem[12165] = 142;
razn_h_mem[12166] = 18;
razn_h_mem[12167] = 148;
razn_h_mem[12168] = 24;
razn_h_mem[12169] = 154;
razn_h_mem[12170] = 30;
razn_h_mem[12171] = 160;
razn_h_mem[12172] = 36;
razn_h_mem[12173] = 166;
razn_h_mem[12174] = 42;
razn_h_mem[12175] = 172;
razn_h_mem[12176] = 48;
razn_h_mem[12177] = 178;
razn_h_mem[12178] = 54;
razn_h_mem[12179] = 184;
razn_h_mem[12180] = 60;
razn_h_mem[12181] = 190;
razn_h_mem[12182] = 66;
razn_h_mem[12183] = 196;
razn_h_mem[12184] = 72;
razn_h_mem[12185] = 202;
razn_h_mem[12186] = 78;
razn_h_mem[12187] = 208;
razn_h_mem[12188] = 84;
razn_h_mem[12189] = 214;
razn_h_mem[12190] = 90;
razn_h_mem[12191] = 220;
razn_h_mem[12192] = 96;
razn_h_mem[12193] = 226;
razn_h_mem[12194] = 102;
razn_h_mem[12195] = 232;
razn_h_mem[12196] = 108;
razn_h_mem[12197] = 238;
razn_h_mem[12198] = 114;
razn_h_mem[12199] = 244;
razn_h_mem[12200] = 120;
razn_h_mem[12201] = 250;
razn_h_mem[12202] = 126;
razn_h_mem[12203] = 2;
razn_h_mem[12204] = 132;
razn_h_mem[12205] = 8;
razn_h_mem[12206] = 138;
razn_h_mem[12207] = 14;
razn_h_mem[12208] = 144;
razn_h_mem[12209] = 20;
razn_h_mem[12210] = 150;
razn_h_mem[12211] = 26;
razn_h_mem[12212] = 156;
razn_h_mem[12213] = 32;
razn_h_mem[12214] = 162;
razn_h_mem[12215] = 38;
razn_h_mem[12216] = 168;
razn_h_mem[12217] = 44;
razn_h_mem[12218] = 174;
razn_h_mem[12219] = 50;
razn_h_mem[12220] = 180;
razn_h_mem[12221] = 56;
razn_h_mem[12222] = 186;
razn_h_mem[12223] = 62;
razn_h_mem[12224] = 192;
razn_h_mem[12225] = 68;
razn_h_mem[12226] = 198;
razn_h_mem[12227] = 74;
razn_h_mem[12228] = 204;
razn_h_mem[12229] = 80;
razn_h_mem[12230] = 210;
razn_h_mem[12231] = 86;
razn_h_mem[12232] = 216;
razn_h_mem[12233] = 92;
razn_h_mem[12234] = 222;
razn_h_mem[12235] = 98;
razn_h_mem[12236] = 228;
razn_h_mem[12237] = 104;
razn_h_mem[12238] = 234;
razn_h_mem[12239] = 110;
razn_h_mem[12240] = 240;
razn_h_mem[12241] = 116;
razn_h_mem[12242] = 246;
razn_h_mem[12243] = 122;
razn_h_mem[12244] = 252;
razn_h_mem[12245] = 128;
razn_h_mem[12246] = 4;
razn_h_mem[12247] = 134;
razn_h_mem[12248] = 10;
razn_h_mem[12249] = 140;
razn_h_mem[12250] = 16;
razn_h_mem[12251] = 146;
razn_h_mem[12252] = 22;
razn_h_mem[12253] = 152;
razn_h_mem[12254] = 28;
razn_h_mem[12255] = 158;
razn_h_mem[12256] = 34;
razn_h_mem[12257] = 164;
razn_h_mem[12258] = 40;
razn_h_mem[12259] = 170;
razn_h_mem[12260] = 46;
razn_h_mem[12261] = 176;
razn_h_mem[12262] = 52;
razn_h_mem[12263] = 182;
razn_h_mem[12264] = 58;
razn_h_mem[12265] = 188;
razn_h_mem[12266] = 64;
razn_h_mem[12267] = 194;
razn_h_mem[12268] = 70;
razn_h_mem[12269] = 200;
razn_h_mem[12270] = 76;
razn_h_mem[12271] = 206;
razn_h_mem[12272] = 82;
razn_h_mem[12273] = 212;
razn_h_mem[12274] = 88;
razn_h_mem[12275] = 218;
razn_h_mem[12276] = 94;
razn_h_mem[12277] = 224;
razn_h_mem[12278] = 100;
razn_h_mem[12279] = 230;
razn_h_mem[12280] = 106;
razn_h_mem[12281] = 236;
razn_h_mem[12282] = 112;
razn_h_mem[12283] = 242;
razn_h_mem[12284] = 118;
razn_h_mem[12285] = 248;
razn_h_mem[12286] = 124;
razn_h_mem[12287] = 255;
razn_h_mem[12288] = 0;
razn_h_mem[12289] = 130;
razn_h_mem[12290] = 6;
razn_h_mem[12291] = 136;
razn_h_mem[12292] = 12;
razn_h_mem[12293] = 142;
razn_h_mem[12294] = 18;
razn_h_mem[12295] = 148;
razn_h_mem[12296] = 24;
razn_h_mem[12297] = 154;
razn_h_mem[12298] = 30;
razn_h_mem[12299] = 160;
razn_h_mem[12300] = 36;
razn_h_mem[12301] = 166;
razn_h_mem[12302] = 42;
razn_h_mem[12303] = 172;
razn_h_mem[12304] = 48;
razn_h_mem[12305] = 178;
razn_h_mem[12306] = 54;
razn_h_mem[12307] = 184;
razn_h_mem[12308] = 60;
razn_h_mem[12309] = 190;
razn_h_mem[12310] = 66;
razn_h_mem[12311] = 196;
razn_h_mem[12312] = 72;
razn_h_mem[12313] = 202;
razn_h_mem[12314] = 78;
razn_h_mem[12315] = 208;
razn_h_mem[12316] = 84;
razn_h_mem[12317] = 214;
razn_h_mem[12318] = 90;
razn_h_mem[12319] = 220;
razn_h_mem[12320] = 96;
razn_h_mem[12321] = 226;
razn_h_mem[12322] = 102;
razn_h_mem[12323] = 232;
razn_h_mem[12324] = 108;
razn_h_mem[12325] = 238;
razn_h_mem[12326] = 114;
razn_h_mem[12327] = 244;
razn_h_mem[12328] = 120;
razn_h_mem[12329] = 250;
razn_h_mem[12330] = 126;
razn_h_mem[12331] = 2;
razn_h_mem[12332] = 132;
razn_h_mem[12333] = 8;
razn_h_mem[12334] = 138;
razn_h_mem[12335] = 14;
razn_h_mem[12336] = 144;
razn_h_mem[12337] = 20;
razn_h_mem[12338] = 150;
razn_h_mem[12339] = 26;
razn_h_mem[12340] = 156;
razn_h_mem[12341] = 32;
razn_h_mem[12342] = 162;
razn_h_mem[12343] = 38;
razn_h_mem[12344] = 168;
razn_h_mem[12345] = 44;
razn_h_mem[12346] = 174;
razn_h_mem[12347] = 50;
razn_h_mem[12348] = 180;
razn_h_mem[12349] = 56;
razn_h_mem[12350] = 186;
razn_h_mem[12351] = 62;
razn_h_mem[12352] = 192;
razn_h_mem[12353] = 68;
razn_h_mem[12354] = 198;
razn_h_mem[12355] = 74;
razn_h_mem[12356] = 204;
razn_h_mem[12357] = 80;
razn_h_mem[12358] = 210;
razn_h_mem[12359] = 86;
razn_h_mem[12360] = 216;
razn_h_mem[12361] = 92;
razn_h_mem[12362] = 222;
razn_h_mem[12363] = 98;
razn_h_mem[12364] = 228;
razn_h_mem[12365] = 104;
razn_h_mem[12366] = 234;
razn_h_mem[12367] = 110;
razn_h_mem[12368] = 240;
razn_h_mem[12369] = 116;
razn_h_mem[12370] = 246;
razn_h_mem[12371] = 122;
razn_h_mem[12372] = 252;
razn_h_mem[12373] = 128;
razn_h_mem[12374] = 4;
razn_h_mem[12375] = 134;
razn_h_mem[12376] = 10;
razn_h_mem[12377] = 140;
razn_h_mem[12378] = 16;
razn_h_mem[12379] = 146;
razn_h_mem[12380] = 22;
razn_h_mem[12381] = 152;
razn_h_mem[12382] = 28;
razn_h_mem[12383] = 158;
razn_h_mem[12384] = 34;
razn_h_mem[12385] = 164;
razn_h_mem[12386] = 40;
razn_h_mem[12387] = 170;
razn_h_mem[12388] = 46;
razn_h_mem[12389] = 176;
razn_h_mem[12390] = 52;
razn_h_mem[12391] = 182;
razn_h_mem[12392] = 58;
razn_h_mem[12393] = 188;
razn_h_mem[12394] = 64;
razn_h_mem[12395] = 194;
razn_h_mem[12396] = 70;
razn_h_mem[12397] = 200;
razn_h_mem[12398] = 76;
razn_h_mem[12399] = 206;
razn_h_mem[12400] = 82;
razn_h_mem[12401] = 212;
razn_h_mem[12402] = 88;
razn_h_mem[12403] = 218;
razn_h_mem[12404] = 94;
razn_h_mem[12405] = 224;
razn_h_mem[12406] = 100;
razn_h_mem[12407] = 230;
razn_h_mem[12408] = 106;
razn_h_mem[12409] = 236;
razn_h_mem[12410] = 112;
razn_h_mem[12411] = 242;
razn_h_mem[12412] = 118;
razn_h_mem[12413] = 248;
razn_h_mem[12414] = 124;
razn_h_mem[12415] = 255;
razn_h_mem[12416] = 0;
razn_h_mem[12417] = 130;
razn_h_mem[12418] = 6;
razn_h_mem[12419] = 136;
razn_h_mem[12420] = 12;
razn_h_mem[12421] = 142;
razn_h_mem[12422] = 18;
razn_h_mem[12423] = 148;
razn_h_mem[12424] = 24;
razn_h_mem[12425] = 154;
razn_h_mem[12426] = 30;
razn_h_mem[12427] = 160;
razn_h_mem[12428] = 36;
razn_h_mem[12429] = 166;
razn_h_mem[12430] = 42;
razn_h_mem[12431] = 172;
razn_h_mem[12432] = 48;
razn_h_mem[12433] = 178;
razn_h_mem[12434] = 54;
razn_h_mem[12435] = 184;
razn_h_mem[12436] = 60;
razn_h_mem[12437] = 190;
razn_h_mem[12438] = 66;
razn_h_mem[12439] = 196;
razn_h_mem[12440] = 72;
razn_h_mem[12441] = 202;
razn_h_mem[12442] = 78;
razn_h_mem[12443] = 208;
razn_h_mem[12444] = 84;
razn_h_mem[12445] = 214;
razn_h_mem[12446] = 90;
razn_h_mem[12447] = 220;
razn_h_mem[12448] = 96;
razn_h_mem[12449] = 226;
razn_h_mem[12450] = 102;
razn_h_mem[12451] = 232;
razn_h_mem[12452] = 108;
razn_h_mem[12453] = 238;
razn_h_mem[12454] = 114;
razn_h_mem[12455] = 244;
razn_h_mem[12456] = 120;
razn_h_mem[12457] = 250;
razn_h_mem[12458] = 126;
razn_h_mem[12459] = 2;
razn_h_mem[12460] = 132;
razn_h_mem[12461] = 8;
razn_h_mem[12462] = 138;
razn_h_mem[12463] = 14;
razn_h_mem[12464] = 144;
razn_h_mem[12465] = 20;
razn_h_mem[12466] = 150;
razn_h_mem[12467] = 26;
razn_h_mem[12468] = 156;
razn_h_mem[12469] = 32;
razn_h_mem[12470] = 162;
razn_h_mem[12471] = 38;
razn_h_mem[12472] = 168;
razn_h_mem[12473] = 44;
razn_h_mem[12474] = 174;
razn_h_mem[12475] = 50;
razn_h_mem[12476] = 180;
razn_h_mem[12477] = 56;
razn_h_mem[12478] = 186;
razn_h_mem[12479] = 62;
razn_h_mem[12480] = 192;
razn_h_mem[12481] = 68;
razn_h_mem[12482] = 198;
razn_h_mem[12483] = 74;
razn_h_mem[12484] = 204;
razn_h_mem[12485] = 80;
razn_h_mem[12486] = 210;
razn_h_mem[12487] = 86;
razn_h_mem[12488] = 216;
razn_h_mem[12489] = 92;
razn_h_mem[12490] = 222;
razn_h_mem[12491] = 98;
razn_h_mem[12492] = 228;
razn_h_mem[12493] = 104;
razn_h_mem[12494] = 234;
razn_h_mem[12495] = 110;
razn_h_mem[12496] = 240;
razn_h_mem[12497] = 116;
razn_h_mem[12498] = 246;
razn_h_mem[12499] = 122;
razn_h_mem[12500] = 252;
razn_h_mem[12501] = 128;
razn_h_mem[12502] = 4;
razn_h_mem[12503] = 134;
razn_h_mem[12504] = 10;
razn_h_mem[12505] = 140;
razn_h_mem[12506] = 16;
razn_h_mem[12507] = 146;
razn_h_mem[12508] = 22;
razn_h_mem[12509] = 152;
razn_h_mem[12510] = 28;
razn_h_mem[12511] = 158;
razn_h_mem[12512] = 34;
razn_h_mem[12513] = 164;
razn_h_mem[12514] = 40;
razn_h_mem[12515] = 170;
razn_h_mem[12516] = 46;
razn_h_mem[12517] = 176;
razn_h_mem[12518] = 52;
razn_h_mem[12519] = 182;
razn_h_mem[12520] = 58;
razn_h_mem[12521] = 188;
razn_h_mem[12522] = 64;
razn_h_mem[12523] = 194;
razn_h_mem[12524] = 70;
razn_h_mem[12525] = 200;
razn_h_mem[12526] = 76;
razn_h_mem[12527] = 206;
razn_h_mem[12528] = 82;
razn_h_mem[12529] = 212;
razn_h_mem[12530] = 88;
razn_h_mem[12531] = 218;
razn_h_mem[12532] = 94;
razn_h_mem[12533] = 224;
razn_h_mem[12534] = 100;
razn_h_mem[12535] = 230;
razn_h_mem[12536] = 106;
razn_h_mem[12537] = 236;
razn_h_mem[12538] = 112;
razn_h_mem[12539] = 242;
razn_h_mem[12540] = 118;
razn_h_mem[12541] = 248;
razn_h_mem[12542] = 124;
razn_h_mem[12543] = 255;
razn_h_mem[12544] = 0;
razn_h_mem[12545] = 130;
razn_h_mem[12546] = 6;
razn_h_mem[12547] = 136;
razn_h_mem[12548] = 12;
razn_h_mem[12549] = 142;
razn_h_mem[12550] = 18;
razn_h_mem[12551] = 148;
razn_h_mem[12552] = 24;
razn_h_mem[12553] = 154;
razn_h_mem[12554] = 30;
razn_h_mem[12555] = 160;
razn_h_mem[12556] = 36;
razn_h_mem[12557] = 166;
razn_h_mem[12558] = 42;
razn_h_mem[12559] = 172;
razn_h_mem[12560] = 48;
razn_h_mem[12561] = 178;
razn_h_mem[12562] = 54;
razn_h_mem[12563] = 184;
razn_h_mem[12564] = 60;
razn_h_mem[12565] = 190;
razn_h_mem[12566] = 66;
razn_h_mem[12567] = 196;
razn_h_mem[12568] = 72;
razn_h_mem[12569] = 202;
razn_h_mem[12570] = 78;
razn_h_mem[12571] = 208;
razn_h_mem[12572] = 84;
razn_h_mem[12573] = 214;
razn_h_mem[12574] = 90;
razn_h_mem[12575] = 220;
razn_h_mem[12576] = 96;
razn_h_mem[12577] = 226;
razn_h_mem[12578] = 102;
razn_h_mem[12579] = 232;
razn_h_mem[12580] = 108;
razn_h_mem[12581] = 238;
razn_h_mem[12582] = 114;
razn_h_mem[12583] = 244;
razn_h_mem[12584] = 120;
razn_h_mem[12585] = 250;
razn_h_mem[12586] = 126;
razn_h_mem[12587] = 2;
razn_h_mem[12588] = 132;
razn_h_mem[12589] = 8;
razn_h_mem[12590] = 138;
razn_h_mem[12591] = 14;
razn_h_mem[12592] = 144;
razn_h_mem[12593] = 20;
razn_h_mem[12594] = 150;
razn_h_mem[12595] = 26;
razn_h_mem[12596] = 156;
razn_h_mem[12597] = 32;
razn_h_mem[12598] = 162;
razn_h_mem[12599] = 38;
razn_h_mem[12600] = 168;
razn_h_mem[12601] = 44;
razn_h_mem[12602] = 174;
razn_h_mem[12603] = 50;
razn_h_mem[12604] = 180;
razn_h_mem[12605] = 56;
razn_h_mem[12606] = 186;
razn_h_mem[12607] = 62;
razn_h_mem[12608] = 192;
razn_h_mem[12609] = 68;
razn_h_mem[12610] = 198;
razn_h_mem[12611] = 74;
razn_h_mem[12612] = 204;
razn_h_mem[12613] = 80;
razn_h_mem[12614] = 210;
razn_h_mem[12615] = 86;
razn_h_mem[12616] = 216;
razn_h_mem[12617] = 92;
razn_h_mem[12618] = 222;
razn_h_mem[12619] = 98;
razn_h_mem[12620] = 228;
razn_h_mem[12621] = 104;
razn_h_mem[12622] = 234;
razn_h_mem[12623] = 110;
razn_h_mem[12624] = 240;
razn_h_mem[12625] = 116;
razn_h_mem[12626] = 246;
razn_h_mem[12627] = 122;
razn_h_mem[12628] = 252;
razn_h_mem[12629] = 128;
razn_h_mem[12630] = 4;
razn_h_mem[12631] = 134;
razn_h_mem[12632] = 10;
razn_h_mem[12633] = 140;
razn_h_mem[12634] = 16;
razn_h_mem[12635] = 146;
razn_h_mem[12636] = 22;
razn_h_mem[12637] = 152;
razn_h_mem[12638] = 28;
razn_h_mem[12639] = 158;
razn_h_mem[12640] = 34;
razn_h_mem[12641] = 164;
razn_h_mem[12642] = 40;
razn_h_mem[12643] = 170;
razn_h_mem[12644] = 46;
razn_h_mem[12645] = 176;
razn_h_mem[12646] = 52;
razn_h_mem[12647] = 182;
razn_h_mem[12648] = 58;
razn_h_mem[12649] = 188;
razn_h_mem[12650] = 64;
razn_h_mem[12651] = 194;
razn_h_mem[12652] = 70;
razn_h_mem[12653] = 200;
razn_h_mem[12654] = 76;
razn_h_mem[12655] = 206;
razn_h_mem[12656] = 82;
razn_h_mem[12657] = 212;
razn_h_mem[12658] = 88;
razn_h_mem[12659] = 218;
razn_h_mem[12660] = 94;
razn_h_mem[12661] = 224;
razn_h_mem[12662] = 100;
razn_h_mem[12663] = 230;
razn_h_mem[12664] = 106;
razn_h_mem[12665] = 236;
razn_h_mem[12666] = 112;
razn_h_mem[12667] = 242;
razn_h_mem[12668] = 118;
razn_h_mem[12669] = 248;
razn_h_mem[12670] = 124;
razn_h_mem[12671] = 255;
razn_h_mem[12672] = 0;
razn_h_mem[12673] = 130;
razn_h_mem[12674] = 6;
razn_h_mem[12675] = 136;
razn_h_mem[12676] = 12;
razn_h_mem[12677] = 142;
razn_h_mem[12678] = 18;
razn_h_mem[12679] = 148;
razn_h_mem[12680] = 24;
razn_h_mem[12681] = 154;
razn_h_mem[12682] = 30;
razn_h_mem[12683] = 160;
razn_h_mem[12684] = 36;
razn_h_mem[12685] = 166;
razn_h_mem[12686] = 42;
razn_h_mem[12687] = 172;
razn_h_mem[12688] = 48;
razn_h_mem[12689] = 178;
razn_h_mem[12690] = 54;
razn_h_mem[12691] = 184;
razn_h_mem[12692] = 60;
razn_h_mem[12693] = 190;
razn_h_mem[12694] = 66;
razn_h_mem[12695] = 196;
razn_h_mem[12696] = 72;
razn_h_mem[12697] = 202;
razn_h_mem[12698] = 78;
razn_h_mem[12699] = 208;
razn_h_mem[12700] = 84;
razn_h_mem[12701] = 214;
razn_h_mem[12702] = 90;
razn_h_mem[12703] = 220;
razn_h_mem[12704] = 96;
razn_h_mem[12705] = 226;
razn_h_mem[12706] = 102;
razn_h_mem[12707] = 232;
razn_h_mem[12708] = 108;
razn_h_mem[12709] = 238;
razn_h_mem[12710] = 114;
razn_h_mem[12711] = 244;
razn_h_mem[12712] = 120;
razn_h_mem[12713] = 250;
razn_h_mem[12714] = 126;
razn_h_mem[12715] = 2;
razn_h_mem[12716] = 132;
razn_h_mem[12717] = 8;
razn_h_mem[12718] = 138;
razn_h_mem[12719] = 14;
razn_h_mem[12720] = 144;
razn_h_mem[12721] = 20;
razn_h_mem[12722] = 150;
razn_h_mem[12723] = 26;
razn_h_mem[12724] = 156;
razn_h_mem[12725] = 32;
razn_h_mem[12726] = 162;
razn_h_mem[12727] = 38;
razn_h_mem[12728] = 168;
razn_h_mem[12729] = 44;
razn_h_mem[12730] = 174;
razn_h_mem[12731] = 50;
razn_h_mem[12732] = 180;
razn_h_mem[12733] = 56;
razn_h_mem[12734] = 186;
razn_h_mem[12735] = 62;
razn_h_mem[12736] = 192;
razn_h_mem[12737] = 68;
razn_h_mem[12738] = 198;
razn_h_mem[12739] = 74;
razn_h_mem[12740] = 204;
razn_h_mem[12741] = 80;
razn_h_mem[12742] = 210;
razn_h_mem[12743] = 86;
razn_h_mem[12744] = 216;
razn_h_mem[12745] = 92;
razn_h_mem[12746] = 222;
razn_h_mem[12747] = 98;
razn_h_mem[12748] = 228;
razn_h_mem[12749] = 104;
razn_h_mem[12750] = 234;
razn_h_mem[12751] = 110;
razn_h_mem[12752] = 240;
razn_h_mem[12753] = 116;
razn_h_mem[12754] = 246;
razn_h_mem[12755] = 122;
razn_h_mem[12756] = 252;
razn_h_mem[12757] = 128;
razn_h_mem[12758] = 4;
razn_h_mem[12759] = 134;
razn_h_mem[12760] = 10;
razn_h_mem[12761] = 140;
razn_h_mem[12762] = 16;
razn_h_mem[12763] = 146;
razn_h_mem[12764] = 22;
razn_h_mem[12765] = 152;
razn_h_mem[12766] = 28;
razn_h_mem[12767] = 158;
razn_h_mem[12768] = 34;
razn_h_mem[12769] = 164;
razn_h_mem[12770] = 40;
razn_h_mem[12771] = 170;
razn_h_mem[12772] = 46;
razn_h_mem[12773] = 176;
razn_h_mem[12774] = 52;
razn_h_mem[12775] = 182;
razn_h_mem[12776] = 58;
razn_h_mem[12777] = 188;
razn_h_mem[12778] = 64;
razn_h_mem[12779] = 194;
razn_h_mem[12780] = 70;
razn_h_mem[12781] = 200;
razn_h_mem[12782] = 76;
razn_h_mem[12783] = 206;
razn_h_mem[12784] = 82;
razn_h_mem[12785] = 212;
razn_h_mem[12786] = 88;
razn_h_mem[12787] = 218;
razn_h_mem[12788] = 94;
razn_h_mem[12789] = 224;
razn_h_mem[12790] = 100;
razn_h_mem[12791] = 230;
razn_h_mem[12792] = 106;
razn_h_mem[12793] = 236;
razn_h_mem[12794] = 112;
razn_h_mem[12795] = 242;
razn_h_mem[12796] = 118;
razn_h_mem[12797] = 248;
razn_h_mem[12798] = 124;
razn_h_mem[12799] = 255;
razn_h_mem[12800] = 0;
razn_h_mem[12801] = 130;
razn_h_mem[12802] = 6;
razn_h_mem[12803] = 136;
razn_h_mem[12804] = 12;
razn_h_mem[12805] = 142;
razn_h_mem[12806] = 18;
razn_h_mem[12807] = 148;
razn_h_mem[12808] = 24;
razn_h_mem[12809] = 154;
razn_h_mem[12810] = 30;
razn_h_mem[12811] = 160;
razn_h_mem[12812] = 36;
razn_h_mem[12813] = 166;
razn_h_mem[12814] = 42;
razn_h_mem[12815] = 172;
razn_h_mem[12816] = 48;
razn_h_mem[12817] = 178;
razn_h_mem[12818] = 54;
razn_h_mem[12819] = 184;
razn_h_mem[12820] = 60;
razn_h_mem[12821] = 190;
razn_h_mem[12822] = 66;
razn_h_mem[12823] = 196;
razn_h_mem[12824] = 72;
razn_h_mem[12825] = 202;
razn_h_mem[12826] = 78;
razn_h_mem[12827] = 208;
razn_h_mem[12828] = 84;
razn_h_mem[12829] = 214;
razn_h_mem[12830] = 90;
razn_h_mem[12831] = 220;
razn_h_mem[12832] = 96;
razn_h_mem[12833] = 226;
razn_h_mem[12834] = 102;
razn_h_mem[12835] = 232;
razn_h_mem[12836] = 108;
razn_h_mem[12837] = 238;
razn_h_mem[12838] = 114;
razn_h_mem[12839] = 244;
razn_h_mem[12840] = 120;
razn_h_mem[12841] = 250;
razn_h_mem[12842] = 126;
razn_h_mem[12843] = 2;
razn_h_mem[12844] = 132;
razn_h_mem[12845] = 8;
razn_h_mem[12846] = 138;
razn_h_mem[12847] = 14;
razn_h_mem[12848] = 144;
razn_h_mem[12849] = 20;
razn_h_mem[12850] = 150;
razn_h_mem[12851] = 26;
razn_h_mem[12852] = 156;
razn_h_mem[12853] = 32;
razn_h_mem[12854] = 162;
razn_h_mem[12855] = 38;
razn_h_mem[12856] = 168;
razn_h_mem[12857] = 44;
razn_h_mem[12858] = 174;
razn_h_mem[12859] = 50;
razn_h_mem[12860] = 180;
razn_h_mem[12861] = 56;
razn_h_mem[12862] = 186;
razn_h_mem[12863] = 62;
razn_h_mem[12864] = 192;
razn_h_mem[12865] = 68;
razn_h_mem[12866] = 198;
razn_h_mem[12867] = 74;
razn_h_mem[12868] = 204;
razn_h_mem[12869] = 80;
razn_h_mem[12870] = 210;
razn_h_mem[12871] = 86;
razn_h_mem[12872] = 216;
razn_h_mem[12873] = 92;
razn_h_mem[12874] = 222;
razn_h_mem[12875] = 98;
razn_h_mem[12876] = 228;
razn_h_mem[12877] = 104;
razn_h_mem[12878] = 234;
razn_h_mem[12879] = 110;
razn_h_mem[12880] = 240;
razn_h_mem[12881] = 116;
razn_h_mem[12882] = 246;
razn_h_mem[12883] = 122;
razn_h_mem[12884] = 252;
razn_h_mem[12885] = 128;
razn_h_mem[12886] = 4;
razn_h_mem[12887] = 134;
razn_h_mem[12888] = 10;
razn_h_mem[12889] = 140;
razn_h_mem[12890] = 16;
razn_h_mem[12891] = 146;
razn_h_mem[12892] = 22;
razn_h_mem[12893] = 152;
razn_h_mem[12894] = 28;
razn_h_mem[12895] = 158;
razn_h_mem[12896] = 34;
razn_h_mem[12897] = 164;
razn_h_mem[12898] = 40;
razn_h_mem[12899] = 170;
razn_h_mem[12900] = 46;
razn_h_mem[12901] = 176;
razn_h_mem[12902] = 52;
razn_h_mem[12903] = 182;
razn_h_mem[12904] = 58;
razn_h_mem[12905] = 188;
razn_h_mem[12906] = 64;
razn_h_mem[12907] = 194;
razn_h_mem[12908] = 70;
razn_h_mem[12909] = 200;
razn_h_mem[12910] = 76;
razn_h_mem[12911] = 206;
razn_h_mem[12912] = 82;
razn_h_mem[12913] = 212;
razn_h_mem[12914] = 88;
razn_h_mem[12915] = 218;
razn_h_mem[12916] = 94;
razn_h_mem[12917] = 224;
razn_h_mem[12918] = 100;
razn_h_mem[12919] = 230;
razn_h_mem[12920] = 106;
razn_h_mem[12921] = 236;
razn_h_mem[12922] = 112;
razn_h_mem[12923] = 242;
razn_h_mem[12924] = 118;
razn_h_mem[12925] = 248;
razn_h_mem[12926] = 124;
razn_h_mem[12927] = 255;
razn_h_mem[12928] = 0;
razn_h_mem[12929] = 130;
razn_h_mem[12930] = 6;
razn_h_mem[12931] = 136;
razn_h_mem[12932] = 12;
razn_h_mem[12933] = 142;
razn_h_mem[12934] = 18;
razn_h_mem[12935] = 148;
razn_h_mem[12936] = 24;
razn_h_mem[12937] = 154;
razn_h_mem[12938] = 30;
razn_h_mem[12939] = 160;
razn_h_mem[12940] = 36;
razn_h_mem[12941] = 166;
razn_h_mem[12942] = 42;
razn_h_mem[12943] = 172;
razn_h_mem[12944] = 48;
razn_h_mem[12945] = 178;
razn_h_mem[12946] = 54;
razn_h_mem[12947] = 184;
razn_h_mem[12948] = 60;
razn_h_mem[12949] = 190;
razn_h_mem[12950] = 66;
razn_h_mem[12951] = 196;
razn_h_mem[12952] = 72;
razn_h_mem[12953] = 202;
razn_h_mem[12954] = 78;
razn_h_mem[12955] = 208;
razn_h_mem[12956] = 84;
razn_h_mem[12957] = 214;
razn_h_mem[12958] = 90;
razn_h_mem[12959] = 220;
razn_h_mem[12960] = 96;
razn_h_mem[12961] = 226;
razn_h_mem[12962] = 102;
razn_h_mem[12963] = 232;
razn_h_mem[12964] = 108;
razn_h_mem[12965] = 238;
razn_h_mem[12966] = 114;
razn_h_mem[12967] = 244;
razn_h_mem[12968] = 120;
razn_h_mem[12969] = 250;
razn_h_mem[12970] = 126;
razn_h_mem[12971] = 2;
razn_h_mem[12972] = 132;
razn_h_mem[12973] = 8;
razn_h_mem[12974] = 138;
razn_h_mem[12975] = 14;
razn_h_mem[12976] = 144;
razn_h_mem[12977] = 20;
razn_h_mem[12978] = 150;
razn_h_mem[12979] = 26;
razn_h_mem[12980] = 156;
razn_h_mem[12981] = 32;
razn_h_mem[12982] = 162;
razn_h_mem[12983] = 38;
razn_h_mem[12984] = 168;
razn_h_mem[12985] = 44;
razn_h_mem[12986] = 174;
razn_h_mem[12987] = 50;
razn_h_mem[12988] = 180;
razn_h_mem[12989] = 56;
razn_h_mem[12990] = 186;
razn_h_mem[12991] = 62;
razn_h_mem[12992] = 192;
razn_h_mem[12993] = 68;
razn_h_mem[12994] = 198;
razn_h_mem[12995] = 74;
razn_h_mem[12996] = 204;
razn_h_mem[12997] = 80;
razn_h_mem[12998] = 210;
razn_h_mem[12999] = 86;
razn_h_mem[13000] = 216;
razn_h_mem[13001] = 92;
razn_h_mem[13002] = 222;
razn_h_mem[13003] = 98;
razn_h_mem[13004] = 228;
razn_h_mem[13005] = 104;
razn_h_mem[13006] = 234;
razn_h_mem[13007] = 110;
razn_h_mem[13008] = 240;
razn_h_mem[13009] = 116;
razn_h_mem[13010] = 246;
razn_h_mem[13011] = 122;
razn_h_mem[13012] = 252;
razn_h_mem[13013] = 128;
razn_h_mem[13014] = 4;
razn_h_mem[13015] = 134;
razn_h_mem[13016] = 10;
razn_h_mem[13017] = 140;
razn_h_mem[13018] = 16;
razn_h_mem[13019] = 146;
razn_h_mem[13020] = 22;
razn_h_mem[13021] = 152;
razn_h_mem[13022] = 28;
razn_h_mem[13023] = 158;
razn_h_mem[13024] = 34;
razn_h_mem[13025] = 164;
razn_h_mem[13026] = 40;
razn_h_mem[13027] = 170;
razn_h_mem[13028] = 46;
razn_h_mem[13029] = 176;
razn_h_mem[13030] = 52;
razn_h_mem[13031] = 182;
razn_h_mem[13032] = 58;
razn_h_mem[13033] = 188;
razn_h_mem[13034] = 64;
razn_h_mem[13035] = 194;
razn_h_mem[13036] = 70;
razn_h_mem[13037] = 200;
razn_h_mem[13038] = 76;
razn_h_mem[13039] = 206;
razn_h_mem[13040] = 82;
razn_h_mem[13041] = 212;
razn_h_mem[13042] = 88;
razn_h_mem[13043] = 218;
razn_h_mem[13044] = 94;
razn_h_mem[13045] = 224;
razn_h_mem[13046] = 100;
razn_h_mem[13047] = 230;
razn_h_mem[13048] = 106;
razn_h_mem[13049] = 236;
razn_h_mem[13050] = 112;
razn_h_mem[13051] = 242;
razn_h_mem[13052] = 118;
razn_h_mem[13053] = 248;
razn_h_mem[13054] = 124;
razn_h_mem[13055] = 255;
razn_h_mem[13056] = 0;
razn_h_mem[13057] = 130;
razn_h_mem[13058] = 6;
razn_h_mem[13059] = 136;
razn_h_mem[13060] = 12;
razn_h_mem[13061] = 142;
razn_h_mem[13062] = 18;
razn_h_mem[13063] = 148;
razn_h_mem[13064] = 24;
razn_h_mem[13065] = 154;
razn_h_mem[13066] = 30;
razn_h_mem[13067] = 160;
razn_h_mem[13068] = 36;
razn_h_mem[13069] = 166;
razn_h_mem[13070] = 42;
razn_h_mem[13071] = 172;
razn_h_mem[13072] = 48;
razn_h_mem[13073] = 178;
razn_h_mem[13074] = 54;
razn_h_mem[13075] = 184;
razn_h_mem[13076] = 60;
razn_h_mem[13077] = 190;
razn_h_mem[13078] = 66;
razn_h_mem[13079] = 196;
razn_h_mem[13080] = 72;
razn_h_mem[13081] = 202;
razn_h_mem[13082] = 78;
razn_h_mem[13083] = 208;
razn_h_mem[13084] = 84;
razn_h_mem[13085] = 214;
razn_h_mem[13086] = 90;
razn_h_mem[13087] = 220;
razn_h_mem[13088] = 96;
razn_h_mem[13089] = 226;
razn_h_mem[13090] = 102;
razn_h_mem[13091] = 232;
razn_h_mem[13092] = 108;
razn_h_mem[13093] = 238;
razn_h_mem[13094] = 114;
razn_h_mem[13095] = 244;
razn_h_mem[13096] = 120;
razn_h_mem[13097] = 250;
razn_h_mem[13098] = 126;
razn_h_mem[13099] = 2;
razn_h_mem[13100] = 132;
razn_h_mem[13101] = 8;
razn_h_mem[13102] = 138;
razn_h_mem[13103] = 14;
razn_h_mem[13104] = 144;
razn_h_mem[13105] = 20;
razn_h_mem[13106] = 150;
razn_h_mem[13107] = 26;
razn_h_mem[13108] = 156;
razn_h_mem[13109] = 32;
razn_h_mem[13110] = 162;
razn_h_mem[13111] = 38;
razn_h_mem[13112] = 168;
razn_h_mem[13113] = 44;
razn_h_mem[13114] = 174;
razn_h_mem[13115] = 50;
razn_h_mem[13116] = 180;
razn_h_mem[13117] = 56;
razn_h_mem[13118] = 186;
razn_h_mem[13119] = 62;
razn_h_mem[13120] = 192;
razn_h_mem[13121] = 68;
razn_h_mem[13122] = 198;
razn_h_mem[13123] = 74;
razn_h_mem[13124] = 204;
razn_h_mem[13125] = 80;
razn_h_mem[13126] = 210;
razn_h_mem[13127] = 86;
razn_h_mem[13128] = 216;
razn_h_mem[13129] = 92;
razn_h_mem[13130] = 222;
razn_h_mem[13131] = 98;
razn_h_mem[13132] = 228;
razn_h_mem[13133] = 104;
razn_h_mem[13134] = 234;
razn_h_mem[13135] = 110;
razn_h_mem[13136] = 240;
razn_h_mem[13137] = 116;
razn_h_mem[13138] = 246;
razn_h_mem[13139] = 122;
razn_h_mem[13140] = 252;
razn_h_mem[13141] = 128;
razn_h_mem[13142] = 4;
razn_h_mem[13143] = 134;
razn_h_mem[13144] = 10;
razn_h_mem[13145] = 140;
razn_h_mem[13146] = 16;
razn_h_mem[13147] = 146;
razn_h_mem[13148] = 22;
razn_h_mem[13149] = 152;
razn_h_mem[13150] = 28;
razn_h_mem[13151] = 158;
razn_h_mem[13152] = 34;
razn_h_mem[13153] = 164;
razn_h_mem[13154] = 40;
razn_h_mem[13155] = 170;
razn_h_mem[13156] = 46;
razn_h_mem[13157] = 176;
razn_h_mem[13158] = 52;
razn_h_mem[13159] = 182;
razn_h_mem[13160] = 58;
razn_h_mem[13161] = 188;
razn_h_mem[13162] = 64;
razn_h_mem[13163] = 194;
razn_h_mem[13164] = 70;
razn_h_mem[13165] = 200;
razn_h_mem[13166] = 76;
razn_h_mem[13167] = 206;
razn_h_mem[13168] = 82;
razn_h_mem[13169] = 212;
razn_h_mem[13170] = 88;
razn_h_mem[13171] = 218;
razn_h_mem[13172] = 94;
razn_h_mem[13173] = 224;
razn_h_mem[13174] = 100;
razn_h_mem[13175] = 230;
razn_h_mem[13176] = 106;
razn_h_mem[13177] = 236;
razn_h_mem[13178] = 112;
razn_h_mem[13179] = 242;
razn_h_mem[13180] = 118;
razn_h_mem[13181] = 248;
razn_h_mem[13182] = 124;
razn_h_mem[13183] = 255;
razn_h_mem[13184] = 0;
razn_h_mem[13185] = 130;
razn_h_mem[13186] = 6;
razn_h_mem[13187] = 136;
razn_h_mem[13188] = 12;
razn_h_mem[13189] = 142;
razn_h_mem[13190] = 18;
razn_h_mem[13191] = 148;
razn_h_mem[13192] = 24;
razn_h_mem[13193] = 154;
razn_h_mem[13194] = 30;
razn_h_mem[13195] = 160;
razn_h_mem[13196] = 36;
razn_h_mem[13197] = 166;
razn_h_mem[13198] = 42;
razn_h_mem[13199] = 172;
razn_h_mem[13200] = 48;
razn_h_mem[13201] = 178;
razn_h_mem[13202] = 54;
razn_h_mem[13203] = 184;
razn_h_mem[13204] = 60;
razn_h_mem[13205] = 190;
razn_h_mem[13206] = 66;
razn_h_mem[13207] = 196;
razn_h_mem[13208] = 72;
razn_h_mem[13209] = 202;
razn_h_mem[13210] = 78;
razn_h_mem[13211] = 208;
razn_h_mem[13212] = 84;
razn_h_mem[13213] = 214;
razn_h_mem[13214] = 90;
razn_h_mem[13215] = 220;
razn_h_mem[13216] = 96;
razn_h_mem[13217] = 226;
razn_h_mem[13218] = 102;
razn_h_mem[13219] = 232;
razn_h_mem[13220] = 108;
razn_h_mem[13221] = 238;
razn_h_mem[13222] = 114;
razn_h_mem[13223] = 244;
razn_h_mem[13224] = 120;
razn_h_mem[13225] = 250;
razn_h_mem[13226] = 126;
razn_h_mem[13227] = 2;
razn_h_mem[13228] = 132;
razn_h_mem[13229] = 8;
razn_h_mem[13230] = 138;
razn_h_mem[13231] = 14;
razn_h_mem[13232] = 144;
razn_h_mem[13233] = 20;
razn_h_mem[13234] = 150;
razn_h_mem[13235] = 26;
razn_h_mem[13236] = 156;
razn_h_mem[13237] = 32;
razn_h_mem[13238] = 162;
razn_h_mem[13239] = 38;
razn_h_mem[13240] = 168;
razn_h_mem[13241] = 44;
razn_h_mem[13242] = 174;
razn_h_mem[13243] = 50;
razn_h_mem[13244] = 180;
razn_h_mem[13245] = 56;
razn_h_mem[13246] = 186;
razn_h_mem[13247] = 62;
razn_h_mem[13248] = 192;
razn_h_mem[13249] = 68;
razn_h_mem[13250] = 198;
razn_h_mem[13251] = 74;
razn_h_mem[13252] = 204;
razn_h_mem[13253] = 80;
razn_h_mem[13254] = 210;
razn_h_mem[13255] = 86;
razn_h_mem[13256] = 216;
razn_h_mem[13257] = 92;
razn_h_mem[13258] = 222;
razn_h_mem[13259] = 98;
razn_h_mem[13260] = 228;
razn_h_mem[13261] = 104;
razn_h_mem[13262] = 234;
razn_h_mem[13263] = 110;
razn_h_mem[13264] = 240;
razn_h_mem[13265] = 116;
razn_h_mem[13266] = 246;
razn_h_mem[13267] = 122;
razn_h_mem[13268] = 252;
razn_h_mem[13269] = 128;
razn_h_mem[13270] = 4;
razn_h_mem[13271] = 134;
razn_h_mem[13272] = 10;
razn_h_mem[13273] = 140;
razn_h_mem[13274] = 16;
razn_h_mem[13275] = 146;
razn_h_mem[13276] = 22;
razn_h_mem[13277] = 152;
razn_h_mem[13278] = 28;
razn_h_mem[13279] = 158;
razn_h_mem[13280] = 34;
razn_h_mem[13281] = 164;
razn_h_mem[13282] = 40;
razn_h_mem[13283] = 170;
razn_h_mem[13284] = 46;
razn_h_mem[13285] = 176;
razn_h_mem[13286] = 52;
razn_h_mem[13287] = 182;
razn_h_mem[13288] = 58;
razn_h_mem[13289] = 188;
razn_h_mem[13290] = 64;
razn_h_mem[13291] = 194;
razn_h_mem[13292] = 70;
razn_h_mem[13293] = 200;
razn_h_mem[13294] = 76;
razn_h_mem[13295] = 206;
razn_h_mem[13296] = 82;
razn_h_mem[13297] = 212;
razn_h_mem[13298] = 88;
razn_h_mem[13299] = 218;
razn_h_mem[13300] = 94;
razn_h_mem[13301] = 224;
razn_h_mem[13302] = 100;
razn_h_mem[13303] = 230;
razn_h_mem[13304] = 106;
razn_h_mem[13305] = 236;
razn_h_mem[13306] = 112;
razn_h_mem[13307] = 242;
razn_h_mem[13308] = 118;
razn_h_mem[13309] = 248;
razn_h_mem[13310] = 124;
razn_h_mem[13311] = 255;
razn_h_mem[13312] = 0;
razn_h_mem[13313] = 130;
razn_h_mem[13314] = 6;
razn_h_mem[13315] = 136;
razn_h_mem[13316] = 12;
razn_h_mem[13317] = 142;
razn_h_mem[13318] = 18;
razn_h_mem[13319] = 148;
razn_h_mem[13320] = 24;
razn_h_mem[13321] = 154;
razn_h_mem[13322] = 30;
razn_h_mem[13323] = 160;
razn_h_mem[13324] = 36;
razn_h_mem[13325] = 166;
razn_h_mem[13326] = 42;
razn_h_mem[13327] = 172;
razn_h_mem[13328] = 48;
razn_h_mem[13329] = 178;
razn_h_mem[13330] = 54;
razn_h_mem[13331] = 184;
razn_h_mem[13332] = 60;
razn_h_mem[13333] = 190;
razn_h_mem[13334] = 66;
razn_h_mem[13335] = 196;
razn_h_mem[13336] = 72;
razn_h_mem[13337] = 202;
razn_h_mem[13338] = 78;
razn_h_mem[13339] = 208;
razn_h_mem[13340] = 84;
razn_h_mem[13341] = 214;
razn_h_mem[13342] = 90;
razn_h_mem[13343] = 220;
razn_h_mem[13344] = 96;
razn_h_mem[13345] = 226;
razn_h_mem[13346] = 102;
razn_h_mem[13347] = 232;
razn_h_mem[13348] = 108;
razn_h_mem[13349] = 238;
razn_h_mem[13350] = 114;
razn_h_mem[13351] = 244;
razn_h_mem[13352] = 120;
razn_h_mem[13353] = 250;
razn_h_mem[13354] = 126;
razn_h_mem[13355] = 2;
razn_h_mem[13356] = 132;
razn_h_mem[13357] = 8;
razn_h_mem[13358] = 138;
razn_h_mem[13359] = 14;
razn_h_mem[13360] = 144;
razn_h_mem[13361] = 20;
razn_h_mem[13362] = 150;
razn_h_mem[13363] = 26;
razn_h_mem[13364] = 156;
razn_h_mem[13365] = 32;
razn_h_mem[13366] = 162;
razn_h_mem[13367] = 38;
razn_h_mem[13368] = 168;
razn_h_mem[13369] = 44;
razn_h_mem[13370] = 174;
razn_h_mem[13371] = 50;
razn_h_mem[13372] = 180;
razn_h_mem[13373] = 56;
razn_h_mem[13374] = 186;
razn_h_mem[13375] = 62;
razn_h_mem[13376] = 192;
razn_h_mem[13377] = 68;
razn_h_mem[13378] = 198;
razn_h_mem[13379] = 74;
razn_h_mem[13380] = 204;
razn_h_mem[13381] = 80;
razn_h_mem[13382] = 210;
razn_h_mem[13383] = 86;
razn_h_mem[13384] = 216;
razn_h_mem[13385] = 92;
razn_h_mem[13386] = 222;
razn_h_mem[13387] = 98;
razn_h_mem[13388] = 228;
razn_h_mem[13389] = 104;
razn_h_mem[13390] = 234;
razn_h_mem[13391] = 110;
razn_h_mem[13392] = 240;
razn_h_mem[13393] = 116;
razn_h_mem[13394] = 246;
razn_h_mem[13395] = 122;
razn_h_mem[13396] = 252;
razn_h_mem[13397] = 128;
razn_h_mem[13398] = 4;
razn_h_mem[13399] = 134;
razn_h_mem[13400] = 10;
razn_h_mem[13401] = 140;
razn_h_mem[13402] = 16;
razn_h_mem[13403] = 146;
razn_h_mem[13404] = 22;
razn_h_mem[13405] = 152;
razn_h_mem[13406] = 28;
razn_h_mem[13407] = 158;
razn_h_mem[13408] = 34;
razn_h_mem[13409] = 164;
razn_h_mem[13410] = 40;
razn_h_mem[13411] = 170;
razn_h_mem[13412] = 46;
razn_h_mem[13413] = 176;
razn_h_mem[13414] = 52;
razn_h_mem[13415] = 182;
razn_h_mem[13416] = 58;
razn_h_mem[13417] = 188;
razn_h_mem[13418] = 64;
razn_h_mem[13419] = 194;
razn_h_mem[13420] = 70;
razn_h_mem[13421] = 200;
razn_h_mem[13422] = 76;
razn_h_mem[13423] = 206;
razn_h_mem[13424] = 82;
razn_h_mem[13425] = 212;
razn_h_mem[13426] = 88;
razn_h_mem[13427] = 218;
razn_h_mem[13428] = 94;
razn_h_mem[13429] = 224;
razn_h_mem[13430] = 100;
razn_h_mem[13431] = 230;
razn_h_mem[13432] = 106;
razn_h_mem[13433] = 236;
razn_h_mem[13434] = 112;
razn_h_mem[13435] = 242;
razn_h_mem[13436] = 118;
razn_h_mem[13437] = 248;
razn_h_mem[13438] = 124;
razn_h_mem[13439] = 255;
razn_h_mem[13440] = 0;
razn_h_mem[13441] = 130;
razn_h_mem[13442] = 6;
razn_h_mem[13443] = 136;
razn_h_mem[13444] = 12;
razn_h_mem[13445] = 142;
razn_h_mem[13446] = 18;
razn_h_mem[13447] = 148;
razn_h_mem[13448] = 24;
razn_h_mem[13449] = 154;
razn_h_mem[13450] = 30;
razn_h_mem[13451] = 160;
razn_h_mem[13452] = 36;
razn_h_mem[13453] = 166;
razn_h_mem[13454] = 42;
razn_h_mem[13455] = 172;
razn_h_mem[13456] = 48;
razn_h_mem[13457] = 178;
razn_h_mem[13458] = 54;
razn_h_mem[13459] = 184;
razn_h_mem[13460] = 60;
razn_h_mem[13461] = 190;
razn_h_mem[13462] = 66;
razn_h_mem[13463] = 196;
razn_h_mem[13464] = 72;
razn_h_mem[13465] = 202;
razn_h_mem[13466] = 78;
razn_h_mem[13467] = 208;
razn_h_mem[13468] = 84;
razn_h_mem[13469] = 214;
razn_h_mem[13470] = 90;
razn_h_mem[13471] = 220;
razn_h_mem[13472] = 96;
razn_h_mem[13473] = 226;
razn_h_mem[13474] = 102;
razn_h_mem[13475] = 232;
razn_h_mem[13476] = 108;
razn_h_mem[13477] = 238;
razn_h_mem[13478] = 114;
razn_h_mem[13479] = 244;
razn_h_mem[13480] = 120;
razn_h_mem[13481] = 250;
razn_h_mem[13482] = 126;
razn_h_mem[13483] = 2;
razn_h_mem[13484] = 132;
razn_h_mem[13485] = 8;
razn_h_mem[13486] = 138;
razn_h_mem[13487] = 14;
razn_h_mem[13488] = 144;
razn_h_mem[13489] = 20;
razn_h_mem[13490] = 150;
razn_h_mem[13491] = 26;
razn_h_mem[13492] = 156;
razn_h_mem[13493] = 32;
razn_h_mem[13494] = 162;
razn_h_mem[13495] = 38;
razn_h_mem[13496] = 168;
razn_h_mem[13497] = 44;
razn_h_mem[13498] = 174;
razn_h_mem[13499] = 50;
razn_h_mem[13500] = 180;
razn_h_mem[13501] = 56;
razn_h_mem[13502] = 186;
razn_h_mem[13503] = 62;
razn_h_mem[13504] = 192;
razn_h_mem[13505] = 68;
razn_h_mem[13506] = 198;
razn_h_mem[13507] = 74;
razn_h_mem[13508] = 204;
razn_h_mem[13509] = 80;
razn_h_mem[13510] = 210;
razn_h_mem[13511] = 86;
razn_h_mem[13512] = 216;
razn_h_mem[13513] = 92;
razn_h_mem[13514] = 222;
razn_h_mem[13515] = 98;
razn_h_mem[13516] = 228;
razn_h_mem[13517] = 104;
razn_h_mem[13518] = 234;
razn_h_mem[13519] = 110;
razn_h_mem[13520] = 240;
razn_h_mem[13521] = 116;
razn_h_mem[13522] = 246;
razn_h_mem[13523] = 122;
razn_h_mem[13524] = 252;
razn_h_mem[13525] = 128;
razn_h_mem[13526] = 4;
razn_h_mem[13527] = 134;
razn_h_mem[13528] = 10;
razn_h_mem[13529] = 140;
razn_h_mem[13530] = 16;
razn_h_mem[13531] = 146;
razn_h_mem[13532] = 22;
razn_h_mem[13533] = 152;
razn_h_mem[13534] = 28;
razn_h_mem[13535] = 158;
razn_h_mem[13536] = 34;
razn_h_mem[13537] = 164;
razn_h_mem[13538] = 40;
razn_h_mem[13539] = 170;
razn_h_mem[13540] = 46;
razn_h_mem[13541] = 176;
razn_h_mem[13542] = 52;
razn_h_mem[13543] = 182;
razn_h_mem[13544] = 58;
razn_h_mem[13545] = 188;
razn_h_mem[13546] = 64;
razn_h_mem[13547] = 194;
razn_h_mem[13548] = 70;
razn_h_mem[13549] = 200;
razn_h_mem[13550] = 76;
razn_h_mem[13551] = 206;
razn_h_mem[13552] = 82;
razn_h_mem[13553] = 212;
razn_h_mem[13554] = 88;
razn_h_mem[13555] = 218;
razn_h_mem[13556] = 94;
razn_h_mem[13557] = 224;
razn_h_mem[13558] = 100;
razn_h_mem[13559] = 230;
razn_h_mem[13560] = 106;
razn_h_mem[13561] = 236;
razn_h_mem[13562] = 112;
razn_h_mem[13563] = 242;
razn_h_mem[13564] = 118;
razn_h_mem[13565] = 248;
razn_h_mem[13566] = 124;
razn_h_mem[13567] = 255;
razn_h_mem[13568] = 0;
razn_h_mem[13569] = 130;
razn_h_mem[13570] = 6;
razn_h_mem[13571] = 136;
razn_h_mem[13572] = 12;
razn_h_mem[13573] = 142;
razn_h_mem[13574] = 18;
razn_h_mem[13575] = 148;
razn_h_mem[13576] = 24;
razn_h_mem[13577] = 154;
razn_h_mem[13578] = 30;
razn_h_mem[13579] = 160;
razn_h_mem[13580] = 36;
razn_h_mem[13581] = 166;
razn_h_mem[13582] = 42;
razn_h_mem[13583] = 172;
razn_h_mem[13584] = 48;
razn_h_mem[13585] = 178;
razn_h_mem[13586] = 54;
razn_h_mem[13587] = 184;
razn_h_mem[13588] = 60;
razn_h_mem[13589] = 190;
razn_h_mem[13590] = 66;
razn_h_mem[13591] = 196;
razn_h_mem[13592] = 72;
razn_h_mem[13593] = 202;
razn_h_mem[13594] = 78;
razn_h_mem[13595] = 208;
razn_h_mem[13596] = 84;
razn_h_mem[13597] = 214;
razn_h_mem[13598] = 90;
razn_h_mem[13599] = 220;
razn_h_mem[13600] = 96;
razn_h_mem[13601] = 226;
razn_h_mem[13602] = 102;
razn_h_mem[13603] = 232;
razn_h_mem[13604] = 108;
razn_h_mem[13605] = 238;
razn_h_mem[13606] = 114;
razn_h_mem[13607] = 244;
razn_h_mem[13608] = 120;
razn_h_mem[13609] = 250;
razn_h_mem[13610] = 126;
razn_h_mem[13611] = 2;
razn_h_mem[13612] = 132;
razn_h_mem[13613] = 8;
razn_h_mem[13614] = 138;
razn_h_mem[13615] = 14;
razn_h_mem[13616] = 144;
razn_h_mem[13617] = 20;
razn_h_mem[13618] = 150;
razn_h_mem[13619] = 26;
razn_h_mem[13620] = 156;
razn_h_mem[13621] = 32;
razn_h_mem[13622] = 162;
razn_h_mem[13623] = 38;
razn_h_mem[13624] = 168;
razn_h_mem[13625] = 44;
razn_h_mem[13626] = 174;
razn_h_mem[13627] = 50;
razn_h_mem[13628] = 180;
razn_h_mem[13629] = 56;
razn_h_mem[13630] = 186;
razn_h_mem[13631] = 62;
razn_h_mem[13632] = 192;
razn_h_mem[13633] = 68;
razn_h_mem[13634] = 198;
razn_h_mem[13635] = 74;
razn_h_mem[13636] = 204;
razn_h_mem[13637] = 80;
razn_h_mem[13638] = 210;
razn_h_mem[13639] = 86;
razn_h_mem[13640] = 216;
razn_h_mem[13641] = 92;
razn_h_mem[13642] = 222;
razn_h_mem[13643] = 98;
razn_h_mem[13644] = 228;
razn_h_mem[13645] = 104;
razn_h_mem[13646] = 234;
razn_h_mem[13647] = 110;
razn_h_mem[13648] = 240;
razn_h_mem[13649] = 116;
razn_h_mem[13650] = 246;
razn_h_mem[13651] = 122;
razn_h_mem[13652] = 252;
razn_h_mem[13653] = 128;
razn_h_mem[13654] = 4;
razn_h_mem[13655] = 134;
razn_h_mem[13656] = 10;
razn_h_mem[13657] = 140;
razn_h_mem[13658] = 16;
razn_h_mem[13659] = 146;
razn_h_mem[13660] = 22;
razn_h_mem[13661] = 152;
razn_h_mem[13662] = 28;
razn_h_mem[13663] = 158;
razn_h_mem[13664] = 34;
razn_h_mem[13665] = 164;
razn_h_mem[13666] = 40;
razn_h_mem[13667] = 170;
razn_h_mem[13668] = 46;
razn_h_mem[13669] = 176;
razn_h_mem[13670] = 52;
razn_h_mem[13671] = 182;
razn_h_mem[13672] = 58;
razn_h_mem[13673] = 188;
razn_h_mem[13674] = 64;
razn_h_mem[13675] = 194;
razn_h_mem[13676] = 70;
razn_h_mem[13677] = 200;
razn_h_mem[13678] = 76;
razn_h_mem[13679] = 206;
razn_h_mem[13680] = 82;
razn_h_mem[13681] = 212;
razn_h_mem[13682] = 88;
razn_h_mem[13683] = 218;
razn_h_mem[13684] = 94;
razn_h_mem[13685] = 224;
razn_h_mem[13686] = 100;
razn_h_mem[13687] = 230;
razn_h_mem[13688] = 106;
razn_h_mem[13689] = 236;
razn_h_mem[13690] = 112;
razn_h_mem[13691] = 242;
razn_h_mem[13692] = 118;
razn_h_mem[13693] = 248;
razn_h_mem[13694] = 124;
razn_h_mem[13695] = 255;
razn_h_mem[13696] = 0;
razn_h_mem[13697] = 130;
razn_h_mem[13698] = 6;
razn_h_mem[13699] = 136;
razn_h_mem[13700] = 12;
razn_h_mem[13701] = 142;
razn_h_mem[13702] = 18;
razn_h_mem[13703] = 148;
razn_h_mem[13704] = 24;
razn_h_mem[13705] = 154;
razn_h_mem[13706] = 30;
razn_h_mem[13707] = 160;
razn_h_mem[13708] = 36;
razn_h_mem[13709] = 166;
razn_h_mem[13710] = 42;
razn_h_mem[13711] = 172;
razn_h_mem[13712] = 48;
razn_h_mem[13713] = 178;
razn_h_mem[13714] = 54;
razn_h_mem[13715] = 184;
razn_h_mem[13716] = 60;
razn_h_mem[13717] = 190;
razn_h_mem[13718] = 66;
razn_h_mem[13719] = 196;
razn_h_mem[13720] = 72;
razn_h_mem[13721] = 202;
razn_h_mem[13722] = 78;
razn_h_mem[13723] = 208;
razn_h_mem[13724] = 84;
razn_h_mem[13725] = 214;
razn_h_mem[13726] = 90;
razn_h_mem[13727] = 220;
razn_h_mem[13728] = 96;
razn_h_mem[13729] = 226;
razn_h_mem[13730] = 102;
razn_h_mem[13731] = 232;
razn_h_mem[13732] = 108;
razn_h_mem[13733] = 238;
razn_h_mem[13734] = 114;
razn_h_mem[13735] = 244;
razn_h_mem[13736] = 120;
razn_h_mem[13737] = 250;
razn_h_mem[13738] = 126;
razn_h_mem[13739] = 2;
razn_h_mem[13740] = 132;
razn_h_mem[13741] = 8;
razn_h_mem[13742] = 138;
razn_h_mem[13743] = 14;
razn_h_mem[13744] = 144;
razn_h_mem[13745] = 20;
razn_h_mem[13746] = 150;
razn_h_mem[13747] = 26;
razn_h_mem[13748] = 156;
razn_h_mem[13749] = 32;
razn_h_mem[13750] = 162;
razn_h_mem[13751] = 38;
razn_h_mem[13752] = 168;
razn_h_mem[13753] = 44;
razn_h_mem[13754] = 174;
razn_h_mem[13755] = 50;
razn_h_mem[13756] = 180;
razn_h_mem[13757] = 56;
razn_h_mem[13758] = 186;
razn_h_mem[13759] = 62;
razn_h_mem[13760] = 192;
razn_h_mem[13761] = 68;
razn_h_mem[13762] = 198;
razn_h_mem[13763] = 74;
razn_h_mem[13764] = 204;
razn_h_mem[13765] = 80;
razn_h_mem[13766] = 210;
razn_h_mem[13767] = 86;
razn_h_mem[13768] = 216;
razn_h_mem[13769] = 92;
razn_h_mem[13770] = 222;
razn_h_mem[13771] = 98;
razn_h_mem[13772] = 228;
razn_h_mem[13773] = 104;
razn_h_mem[13774] = 234;
razn_h_mem[13775] = 110;
razn_h_mem[13776] = 240;
razn_h_mem[13777] = 116;
razn_h_mem[13778] = 246;
razn_h_mem[13779] = 122;
razn_h_mem[13780] = 252;
razn_h_mem[13781] = 128;
razn_h_mem[13782] = 4;
razn_h_mem[13783] = 134;
razn_h_mem[13784] = 10;
razn_h_mem[13785] = 140;
razn_h_mem[13786] = 16;
razn_h_mem[13787] = 146;
razn_h_mem[13788] = 22;
razn_h_mem[13789] = 152;
razn_h_mem[13790] = 28;
razn_h_mem[13791] = 158;
razn_h_mem[13792] = 34;
razn_h_mem[13793] = 164;
razn_h_mem[13794] = 40;
razn_h_mem[13795] = 170;
razn_h_mem[13796] = 46;
razn_h_mem[13797] = 176;
razn_h_mem[13798] = 52;
razn_h_mem[13799] = 182;
razn_h_mem[13800] = 58;
razn_h_mem[13801] = 188;
razn_h_mem[13802] = 64;
razn_h_mem[13803] = 194;
razn_h_mem[13804] = 70;
razn_h_mem[13805] = 200;
razn_h_mem[13806] = 76;
razn_h_mem[13807] = 206;
razn_h_mem[13808] = 82;
razn_h_mem[13809] = 212;
razn_h_mem[13810] = 88;
razn_h_mem[13811] = 218;
razn_h_mem[13812] = 94;
razn_h_mem[13813] = 224;
razn_h_mem[13814] = 100;
razn_h_mem[13815] = 230;
razn_h_mem[13816] = 106;
razn_h_mem[13817] = 236;
razn_h_mem[13818] = 112;
razn_h_mem[13819] = 242;
razn_h_mem[13820] = 118;
razn_h_mem[13821] = 248;
razn_h_mem[13822] = 124;
razn_h_mem[13823] = 255;
razn_h_mem[13824] = 0;
razn_h_mem[13825] = 130;
razn_h_mem[13826] = 6;
razn_h_mem[13827] = 136;
razn_h_mem[13828] = 12;
razn_h_mem[13829] = 142;
razn_h_mem[13830] = 18;
razn_h_mem[13831] = 148;
razn_h_mem[13832] = 24;
razn_h_mem[13833] = 154;
razn_h_mem[13834] = 30;
razn_h_mem[13835] = 160;
razn_h_mem[13836] = 36;
razn_h_mem[13837] = 166;
razn_h_mem[13838] = 42;
razn_h_mem[13839] = 172;
razn_h_mem[13840] = 48;
razn_h_mem[13841] = 178;
razn_h_mem[13842] = 54;
razn_h_mem[13843] = 184;
razn_h_mem[13844] = 60;
razn_h_mem[13845] = 190;
razn_h_mem[13846] = 66;
razn_h_mem[13847] = 196;
razn_h_mem[13848] = 72;
razn_h_mem[13849] = 202;
razn_h_mem[13850] = 78;
razn_h_mem[13851] = 208;
razn_h_mem[13852] = 84;
razn_h_mem[13853] = 214;
razn_h_mem[13854] = 90;
razn_h_mem[13855] = 220;
razn_h_mem[13856] = 96;
razn_h_mem[13857] = 226;
razn_h_mem[13858] = 102;
razn_h_mem[13859] = 232;
razn_h_mem[13860] = 108;
razn_h_mem[13861] = 238;
razn_h_mem[13862] = 114;
razn_h_mem[13863] = 244;
razn_h_mem[13864] = 120;
razn_h_mem[13865] = 250;
razn_h_mem[13866] = 126;
razn_h_mem[13867] = 2;
razn_h_mem[13868] = 132;
razn_h_mem[13869] = 8;
razn_h_mem[13870] = 138;
razn_h_mem[13871] = 14;
razn_h_mem[13872] = 144;
razn_h_mem[13873] = 20;
razn_h_mem[13874] = 150;
razn_h_mem[13875] = 26;
razn_h_mem[13876] = 156;
razn_h_mem[13877] = 32;
razn_h_mem[13878] = 162;
razn_h_mem[13879] = 38;
razn_h_mem[13880] = 168;
razn_h_mem[13881] = 44;
razn_h_mem[13882] = 174;
razn_h_mem[13883] = 50;
razn_h_mem[13884] = 180;
razn_h_mem[13885] = 56;
razn_h_mem[13886] = 186;
razn_h_mem[13887] = 62;
razn_h_mem[13888] = 192;
razn_h_mem[13889] = 68;
razn_h_mem[13890] = 198;
razn_h_mem[13891] = 74;
razn_h_mem[13892] = 204;
razn_h_mem[13893] = 80;
razn_h_mem[13894] = 210;
razn_h_mem[13895] = 86;
razn_h_mem[13896] = 216;
razn_h_mem[13897] = 92;
razn_h_mem[13898] = 222;
razn_h_mem[13899] = 98;
razn_h_mem[13900] = 228;
razn_h_mem[13901] = 104;
razn_h_mem[13902] = 234;
razn_h_mem[13903] = 110;
razn_h_mem[13904] = 240;
razn_h_mem[13905] = 116;
razn_h_mem[13906] = 246;
razn_h_mem[13907] = 122;
razn_h_mem[13908] = 252;
razn_h_mem[13909] = 128;
razn_h_mem[13910] = 4;
razn_h_mem[13911] = 134;
razn_h_mem[13912] = 10;
razn_h_mem[13913] = 140;
razn_h_mem[13914] = 16;
razn_h_mem[13915] = 146;
razn_h_mem[13916] = 22;
razn_h_mem[13917] = 152;
razn_h_mem[13918] = 28;
razn_h_mem[13919] = 158;
razn_h_mem[13920] = 34;
razn_h_mem[13921] = 164;
razn_h_mem[13922] = 40;
razn_h_mem[13923] = 170;
razn_h_mem[13924] = 46;
razn_h_mem[13925] = 176;
razn_h_mem[13926] = 52;
razn_h_mem[13927] = 182;
razn_h_mem[13928] = 58;
razn_h_mem[13929] = 188;
razn_h_mem[13930] = 64;
razn_h_mem[13931] = 194;
razn_h_mem[13932] = 70;
razn_h_mem[13933] = 200;
razn_h_mem[13934] = 76;
razn_h_mem[13935] = 206;
razn_h_mem[13936] = 82;
razn_h_mem[13937] = 212;
razn_h_mem[13938] = 88;
razn_h_mem[13939] = 218;
razn_h_mem[13940] = 94;
razn_h_mem[13941] = 224;
razn_h_mem[13942] = 100;
razn_h_mem[13943] = 230;
razn_h_mem[13944] = 106;
razn_h_mem[13945] = 236;
razn_h_mem[13946] = 112;
razn_h_mem[13947] = 242;
razn_h_mem[13948] = 118;
razn_h_mem[13949] = 248;
razn_h_mem[13950] = 124;
razn_h_mem[13951] = 255;
razn_h_mem[13952] = 0;
razn_h_mem[13953] = 130;
razn_h_mem[13954] = 6;
razn_h_mem[13955] = 136;
razn_h_mem[13956] = 12;
razn_h_mem[13957] = 142;
razn_h_mem[13958] = 18;
razn_h_mem[13959] = 148;
razn_h_mem[13960] = 24;
razn_h_mem[13961] = 154;
razn_h_mem[13962] = 30;
razn_h_mem[13963] = 160;
razn_h_mem[13964] = 36;
razn_h_mem[13965] = 166;
razn_h_mem[13966] = 42;
razn_h_mem[13967] = 172;
razn_h_mem[13968] = 48;
razn_h_mem[13969] = 178;
razn_h_mem[13970] = 54;
razn_h_mem[13971] = 184;
razn_h_mem[13972] = 60;
razn_h_mem[13973] = 190;
razn_h_mem[13974] = 66;
razn_h_mem[13975] = 196;
razn_h_mem[13976] = 72;
razn_h_mem[13977] = 202;
razn_h_mem[13978] = 78;
razn_h_mem[13979] = 208;
razn_h_mem[13980] = 84;
razn_h_mem[13981] = 214;
razn_h_mem[13982] = 90;
razn_h_mem[13983] = 220;
razn_h_mem[13984] = 96;
razn_h_mem[13985] = 226;
razn_h_mem[13986] = 102;
razn_h_mem[13987] = 232;
razn_h_mem[13988] = 108;
razn_h_mem[13989] = 238;
razn_h_mem[13990] = 114;
razn_h_mem[13991] = 244;
razn_h_mem[13992] = 120;
razn_h_mem[13993] = 250;
razn_h_mem[13994] = 126;
razn_h_mem[13995] = 2;
razn_h_mem[13996] = 132;
razn_h_mem[13997] = 8;
razn_h_mem[13998] = 138;
razn_h_mem[13999] = 14;
razn_h_mem[14000] = 144;
razn_h_mem[14001] = 20;
razn_h_mem[14002] = 150;
razn_h_mem[14003] = 26;
razn_h_mem[14004] = 156;
razn_h_mem[14005] = 32;
razn_h_mem[14006] = 162;
razn_h_mem[14007] = 38;
razn_h_mem[14008] = 168;
razn_h_mem[14009] = 44;
razn_h_mem[14010] = 174;
razn_h_mem[14011] = 50;
razn_h_mem[14012] = 180;
razn_h_mem[14013] = 56;
razn_h_mem[14014] = 186;
razn_h_mem[14015] = 62;
razn_h_mem[14016] = 192;
razn_h_mem[14017] = 68;
razn_h_mem[14018] = 198;
razn_h_mem[14019] = 74;
razn_h_mem[14020] = 204;
razn_h_mem[14021] = 80;
razn_h_mem[14022] = 210;
razn_h_mem[14023] = 86;
razn_h_mem[14024] = 216;
razn_h_mem[14025] = 92;
razn_h_mem[14026] = 222;
razn_h_mem[14027] = 98;
razn_h_mem[14028] = 228;
razn_h_mem[14029] = 104;
razn_h_mem[14030] = 234;
razn_h_mem[14031] = 110;
razn_h_mem[14032] = 240;
razn_h_mem[14033] = 116;
razn_h_mem[14034] = 246;
razn_h_mem[14035] = 122;
razn_h_mem[14036] = 252;
razn_h_mem[14037] = 128;
razn_h_mem[14038] = 4;
razn_h_mem[14039] = 134;
razn_h_mem[14040] = 10;
razn_h_mem[14041] = 140;
razn_h_mem[14042] = 16;
razn_h_mem[14043] = 146;
razn_h_mem[14044] = 22;
razn_h_mem[14045] = 152;
razn_h_mem[14046] = 28;
razn_h_mem[14047] = 158;
razn_h_mem[14048] = 34;
razn_h_mem[14049] = 164;
razn_h_mem[14050] = 40;
razn_h_mem[14051] = 170;
razn_h_mem[14052] = 46;
razn_h_mem[14053] = 176;
razn_h_mem[14054] = 52;
razn_h_mem[14055] = 182;
razn_h_mem[14056] = 58;
razn_h_mem[14057] = 188;
razn_h_mem[14058] = 64;
razn_h_mem[14059] = 194;
razn_h_mem[14060] = 70;
razn_h_mem[14061] = 200;
razn_h_mem[14062] = 76;
razn_h_mem[14063] = 206;
razn_h_mem[14064] = 82;
razn_h_mem[14065] = 212;
razn_h_mem[14066] = 88;
razn_h_mem[14067] = 218;
razn_h_mem[14068] = 94;
razn_h_mem[14069] = 224;
razn_h_mem[14070] = 100;
razn_h_mem[14071] = 230;
razn_h_mem[14072] = 106;
razn_h_mem[14073] = 236;
razn_h_mem[14074] = 112;
razn_h_mem[14075] = 242;
razn_h_mem[14076] = 118;
razn_h_mem[14077] = 248;
razn_h_mem[14078] = 124;
razn_h_mem[14079] = 255;
razn_h_mem[14080] = 0;
razn_h_mem[14081] = 130;
razn_h_mem[14082] = 6;
razn_h_mem[14083] = 136;
razn_h_mem[14084] = 12;
razn_h_mem[14085] = 142;
razn_h_mem[14086] = 18;
razn_h_mem[14087] = 148;
razn_h_mem[14088] = 24;
razn_h_mem[14089] = 154;
razn_h_mem[14090] = 30;
razn_h_mem[14091] = 160;
razn_h_mem[14092] = 36;
razn_h_mem[14093] = 166;
razn_h_mem[14094] = 42;
razn_h_mem[14095] = 172;
razn_h_mem[14096] = 48;
razn_h_mem[14097] = 178;
razn_h_mem[14098] = 54;
razn_h_mem[14099] = 184;
razn_h_mem[14100] = 60;
razn_h_mem[14101] = 190;
razn_h_mem[14102] = 66;
razn_h_mem[14103] = 196;
razn_h_mem[14104] = 72;
razn_h_mem[14105] = 202;
razn_h_mem[14106] = 78;
razn_h_mem[14107] = 208;
razn_h_mem[14108] = 84;
razn_h_mem[14109] = 214;
razn_h_mem[14110] = 90;
razn_h_mem[14111] = 220;
razn_h_mem[14112] = 96;
razn_h_mem[14113] = 226;
razn_h_mem[14114] = 102;
razn_h_mem[14115] = 232;
razn_h_mem[14116] = 108;
razn_h_mem[14117] = 238;
razn_h_mem[14118] = 114;
razn_h_mem[14119] = 244;
razn_h_mem[14120] = 120;
razn_h_mem[14121] = 250;
razn_h_mem[14122] = 126;
razn_h_mem[14123] = 2;
razn_h_mem[14124] = 132;
razn_h_mem[14125] = 8;
razn_h_mem[14126] = 138;
razn_h_mem[14127] = 14;
razn_h_mem[14128] = 144;
razn_h_mem[14129] = 20;
razn_h_mem[14130] = 150;
razn_h_mem[14131] = 26;
razn_h_mem[14132] = 156;
razn_h_mem[14133] = 32;
razn_h_mem[14134] = 162;
razn_h_mem[14135] = 38;
razn_h_mem[14136] = 168;
razn_h_mem[14137] = 44;
razn_h_mem[14138] = 174;
razn_h_mem[14139] = 50;
razn_h_mem[14140] = 180;
razn_h_mem[14141] = 56;
razn_h_mem[14142] = 186;
razn_h_mem[14143] = 62;
razn_h_mem[14144] = 192;
razn_h_mem[14145] = 68;
razn_h_mem[14146] = 198;
razn_h_mem[14147] = 74;
razn_h_mem[14148] = 204;
razn_h_mem[14149] = 80;
razn_h_mem[14150] = 210;
razn_h_mem[14151] = 86;
razn_h_mem[14152] = 216;
razn_h_mem[14153] = 92;
razn_h_mem[14154] = 222;
razn_h_mem[14155] = 98;
razn_h_mem[14156] = 228;
razn_h_mem[14157] = 104;
razn_h_mem[14158] = 234;
razn_h_mem[14159] = 110;
razn_h_mem[14160] = 240;
razn_h_mem[14161] = 116;
razn_h_mem[14162] = 246;
razn_h_mem[14163] = 122;
razn_h_mem[14164] = 252;
razn_h_mem[14165] = 128;
razn_h_mem[14166] = 4;
razn_h_mem[14167] = 134;
razn_h_mem[14168] = 10;
razn_h_mem[14169] = 140;
razn_h_mem[14170] = 16;
razn_h_mem[14171] = 146;
razn_h_mem[14172] = 22;
razn_h_mem[14173] = 152;
razn_h_mem[14174] = 28;
razn_h_mem[14175] = 158;
razn_h_mem[14176] = 34;
razn_h_mem[14177] = 164;
razn_h_mem[14178] = 40;
razn_h_mem[14179] = 170;
razn_h_mem[14180] = 46;
razn_h_mem[14181] = 176;
razn_h_mem[14182] = 52;
razn_h_mem[14183] = 182;
razn_h_mem[14184] = 58;
razn_h_mem[14185] = 188;
razn_h_mem[14186] = 64;
razn_h_mem[14187] = 194;
razn_h_mem[14188] = 70;
razn_h_mem[14189] = 200;
razn_h_mem[14190] = 76;
razn_h_mem[14191] = 206;
razn_h_mem[14192] = 82;
razn_h_mem[14193] = 212;
razn_h_mem[14194] = 88;
razn_h_mem[14195] = 218;
razn_h_mem[14196] = 94;
razn_h_mem[14197] = 224;
razn_h_mem[14198] = 100;
razn_h_mem[14199] = 230;
razn_h_mem[14200] = 106;
razn_h_mem[14201] = 236;
razn_h_mem[14202] = 112;
razn_h_mem[14203] = 242;
razn_h_mem[14204] = 118;
razn_h_mem[14205] = 248;
razn_h_mem[14206] = 124;
razn_h_mem[14207] = 255;
razn_h_mem[14208] = 0;
razn_h_mem[14209] = 130;
razn_h_mem[14210] = 6;
razn_h_mem[14211] = 136;
razn_h_mem[14212] = 12;
razn_h_mem[14213] = 142;
razn_h_mem[14214] = 18;
razn_h_mem[14215] = 148;
razn_h_mem[14216] = 24;
razn_h_mem[14217] = 154;
razn_h_mem[14218] = 30;
razn_h_mem[14219] = 160;
razn_h_mem[14220] = 36;
razn_h_mem[14221] = 166;
razn_h_mem[14222] = 42;
razn_h_mem[14223] = 172;
razn_h_mem[14224] = 48;
razn_h_mem[14225] = 178;
razn_h_mem[14226] = 54;
razn_h_mem[14227] = 184;
razn_h_mem[14228] = 60;
razn_h_mem[14229] = 190;
razn_h_mem[14230] = 66;
razn_h_mem[14231] = 196;
razn_h_mem[14232] = 72;
razn_h_mem[14233] = 202;
razn_h_mem[14234] = 78;
razn_h_mem[14235] = 208;
razn_h_mem[14236] = 84;
razn_h_mem[14237] = 214;
razn_h_mem[14238] = 90;
razn_h_mem[14239] = 220;
razn_h_mem[14240] = 96;
razn_h_mem[14241] = 226;
razn_h_mem[14242] = 102;
razn_h_mem[14243] = 232;
razn_h_mem[14244] = 108;
razn_h_mem[14245] = 238;
razn_h_mem[14246] = 114;
razn_h_mem[14247] = 244;
razn_h_mem[14248] = 120;
razn_h_mem[14249] = 250;
razn_h_mem[14250] = 126;
razn_h_mem[14251] = 2;
razn_h_mem[14252] = 132;
razn_h_mem[14253] = 8;
razn_h_mem[14254] = 138;
razn_h_mem[14255] = 14;
razn_h_mem[14256] = 144;
razn_h_mem[14257] = 20;
razn_h_mem[14258] = 150;
razn_h_mem[14259] = 26;
razn_h_mem[14260] = 156;
razn_h_mem[14261] = 32;
razn_h_mem[14262] = 162;
razn_h_mem[14263] = 38;
razn_h_mem[14264] = 168;
razn_h_mem[14265] = 44;
razn_h_mem[14266] = 174;
razn_h_mem[14267] = 50;
razn_h_mem[14268] = 180;
razn_h_mem[14269] = 56;
razn_h_mem[14270] = 186;
razn_h_mem[14271] = 62;
razn_h_mem[14272] = 192;
razn_h_mem[14273] = 68;
razn_h_mem[14274] = 198;
razn_h_mem[14275] = 74;
razn_h_mem[14276] = 204;
razn_h_mem[14277] = 80;
razn_h_mem[14278] = 210;
razn_h_mem[14279] = 86;
razn_h_mem[14280] = 216;
razn_h_mem[14281] = 92;
razn_h_mem[14282] = 222;
razn_h_mem[14283] = 98;
razn_h_mem[14284] = 228;
razn_h_mem[14285] = 104;
razn_h_mem[14286] = 234;
razn_h_mem[14287] = 110;
razn_h_mem[14288] = 240;
razn_h_mem[14289] = 116;
razn_h_mem[14290] = 246;
razn_h_mem[14291] = 122;
razn_h_mem[14292] = 252;
razn_h_mem[14293] = 128;
razn_h_mem[14294] = 4;
razn_h_mem[14295] = 134;
razn_h_mem[14296] = 10;
razn_h_mem[14297] = 140;
razn_h_mem[14298] = 16;
razn_h_mem[14299] = 146;
razn_h_mem[14300] = 22;
razn_h_mem[14301] = 152;
razn_h_mem[14302] = 28;
razn_h_mem[14303] = 158;
razn_h_mem[14304] = 34;
razn_h_mem[14305] = 164;
razn_h_mem[14306] = 40;
razn_h_mem[14307] = 170;
razn_h_mem[14308] = 46;
razn_h_mem[14309] = 176;
razn_h_mem[14310] = 52;
razn_h_mem[14311] = 182;
razn_h_mem[14312] = 58;
razn_h_mem[14313] = 188;
razn_h_mem[14314] = 64;
razn_h_mem[14315] = 194;
razn_h_mem[14316] = 70;
razn_h_mem[14317] = 200;
razn_h_mem[14318] = 76;
razn_h_mem[14319] = 206;
razn_h_mem[14320] = 82;
razn_h_mem[14321] = 212;
razn_h_mem[14322] = 88;
razn_h_mem[14323] = 218;
razn_h_mem[14324] = 94;
razn_h_mem[14325] = 224;
razn_h_mem[14326] = 100;
razn_h_mem[14327] = 230;
razn_h_mem[14328] = 106;
razn_h_mem[14329] = 236;
razn_h_mem[14330] = 112;
razn_h_mem[14331] = 242;
razn_h_mem[14332] = 118;
razn_h_mem[14333] = 248;
razn_h_mem[14334] = 124;
razn_h_mem[14335] = 255;
razn_h_mem[14336] = 0;
razn_h_mem[14337] = 130;
razn_h_mem[14338] = 6;
razn_h_mem[14339] = 136;
razn_h_mem[14340] = 12;
razn_h_mem[14341] = 142;
razn_h_mem[14342] = 18;
razn_h_mem[14343] = 148;
razn_h_mem[14344] = 24;
razn_h_mem[14345] = 154;
razn_h_mem[14346] = 30;
razn_h_mem[14347] = 160;
razn_h_mem[14348] = 36;
razn_h_mem[14349] = 166;
razn_h_mem[14350] = 42;
razn_h_mem[14351] = 172;
razn_h_mem[14352] = 48;
razn_h_mem[14353] = 178;
razn_h_mem[14354] = 54;
razn_h_mem[14355] = 184;
razn_h_mem[14356] = 60;
razn_h_mem[14357] = 190;
razn_h_mem[14358] = 66;
razn_h_mem[14359] = 196;
razn_h_mem[14360] = 72;
razn_h_mem[14361] = 202;
razn_h_mem[14362] = 78;
razn_h_mem[14363] = 208;
razn_h_mem[14364] = 84;
razn_h_mem[14365] = 214;
razn_h_mem[14366] = 90;
razn_h_mem[14367] = 220;
razn_h_mem[14368] = 96;
razn_h_mem[14369] = 226;
razn_h_mem[14370] = 102;
razn_h_mem[14371] = 232;
razn_h_mem[14372] = 108;
razn_h_mem[14373] = 238;
razn_h_mem[14374] = 114;
razn_h_mem[14375] = 244;
razn_h_mem[14376] = 120;
razn_h_mem[14377] = 250;
razn_h_mem[14378] = 126;
razn_h_mem[14379] = 2;
razn_h_mem[14380] = 132;
razn_h_mem[14381] = 8;
razn_h_mem[14382] = 138;
razn_h_mem[14383] = 14;
razn_h_mem[14384] = 144;
razn_h_mem[14385] = 20;
razn_h_mem[14386] = 150;
razn_h_mem[14387] = 26;
razn_h_mem[14388] = 156;
razn_h_mem[14389] = 32;
razn_h_mem[14390] = 162;
razn_h_mem[14391] = 38;
razn_h_mem[14392] = 168;
razn_h_mem[14393] = 44;
razn_h_mem[14394] = 174;
razn_h_mem[14395] = 50;
razn_h_mem[14396] = 180;
razn_h_mem[14397] = 56;
razn_h_mem[14398] = 186;
razn_h_mem[14399] = 62;
razn_h_mem[14400] = 192;
razn_h_mem[14401] = 68;
razn_h_mem[14402] = 198;
razn_h_mem[14403] = 74;
razn_h_mem[14404] = 204;
razn_h_mem[14405] = 80;
razn_h_mem[14406] = 210;
razn_h_mem[14407] = 86;
razn_h_mem[14408] = 216;
razn_h_mem[14409] = 92;
razn_h_mem[14410] = 222;
razn_h_mem[14411] = 98;
razn_h_mem[14412] = 228;
razn_h_mem[14413] = 104;
razn_h_mem[14414] = 234;
razn_h_mem[14415] = 110;
razn_h_mem[14416] = 240;
razn_h_mem[14417] = 116;
razn_h_mem[14418] = 246;
razn_h_mem[14419] = 122;
razn_h_mem[14420] = 252;
razn_h_mem[14421] = 128;
razn_h_mem[14422] = 4;
razn_h_mem[14423] = 134;
razn_h_mem[14424] = 10;
razn_h_mem[14425] = 140;
razn_h_mem[14426] = 16;
razn_h_mem[14427] = 146;
razn_h_mem[14428] = 22;
razn_h_mem[14429] = 152;
razn_h_mem[14430] = 28;
razn_h_mem[14431] = 158;
razn_h_mem[14432] = 34;
razn_h_mem[14433] = 164;
razn_h_mem[14434] = 40;
razn_h_mem[14435] = 170;
razn_h_mem[14436] = 46;
razn_h_mem[14437] = 176;
razn_h_mem[14438] = 52;
razn_h_mem[14439] = 182;
razn_h_mem[14440] = 58;
razn_h_mem[14441] = 188;
razn_h_mem[14442] = 64;
razn_h_mem[14443] = 194;
razn_h_mem[14444] = 70;
razn_h_mem[14445] = 200;
razn_h_mem[14446] = 76;
razn_h_mem[14447] = 206;
razn_h_mem[14448] = 82;
razn_h_mem[14449] = 212;
razn_h_mem[14450] = 88;
razn_h_mem[14451] = 218;
razn_h_mem[14452] = 94;
razn_h_mem[14453] = 224;
razn_h_mem[14454] = 100;
razn_h_mem[14455] = 230;
razn_h_mem[14456] = 106;
razn_h_mem[14457] = 236;
razn_h_mem[14458] = 112;
razn_h_mem[14459] = 242;
razn_h_mem[14460] = 118;
razn_h_mem[14461] = 248;
razn_h_mem[14462] = 124;
razn_h_mem[14463] = 255;
razn_h_mem[14464] = 0;
razn_h_mem[14465] = 130;
razn_h_mem[14466] = 6;
razn_h_mem[14467] = 136;
razn_h_mem[14468] = 12;
razn_h_mem[14469] = 142;
razn_h_mem[14470] = 18;
razn_h_mem[14471] = 148;
razn_h_mem[14472] = 24;
razn_h_mem[14473] = 154;
razn_h_mem[14474] = 30;
razn_h_mem[14475] = 160;
razn_h_mem[14476] = 36;
razn_h_mem[14477] = 166;
razn_h_mem[14478] = 42;
razn_h_mem[14479] = 172;
razn_h_mem[14480] = 48;
razn_h_mem[14481] = 178;
razn_h_mem[14482] = 54;
razn_h_mem[14483] = 184;
razn_h_mem[14484] = 60;
razn_h_mem[14485] = 190;
razn_h_mem[14486] = 66;
razn_h_mem[14487] = 196;
razn_h_mem[14488] = 72;
razn_h_mem[14489] = 202;
razn_h_mem[14490] = 78;
razn_h_mem[14491] = 208;
razn_h_mem[14492] = 84;
razn_h_mem[14493] = 214;
razn_h_mem[14494] = 90;
razn_h_mem[14495] = 220;
razn_h_mem[14496] = 96;
razn_h_mem[14497] = 226;
razn_h_mem[14498] = 102;
razn_h_mem[14499] = 232;
razn_h_mem[14500] = 108;
razn_h_mem[14501] = 238;
razn_h_mem[14502] = 114;
razn_h_mem[14503] = 244;
razn_h_mem[14504] = 120;
razn_h_mem[14505] = 250;
razn_h_mem[14506] = 126;
razn_h_mem[14507] = 2;
razn_h_mem[14508] = 132;
razn_h_mem[14509] = 8;
razn_h_mem[14510] = 138;
razn_h_mem[14511] = 14;
razn_h_mem[14512] = 144;
razn_h_mem[14513] = 20;
razn_h_mem[14514] = 150;
razn_h_mem[14515] = 26;
razn_h_mem[14516] = 156;
razn_h_mem[14517] = 32;
razn_h_mem[14518] = 162;
razn_h_mem[14519] = 38;
razn_h_mem[14520] = 168;
razn_h_mem[14521] = 44;
razn_h_mem[14522] = 174;
razn_h_mem[14523] = 50;
razn_h_mem[14524] = 180;
razn_h_mem[14525] = 56;
razn_h_mem[14526] = 186;
razn_h_mem[14527] = 62;
razn_h_mem[14528] = 192;
razn_h_mem[14529] = 68;
razn_h_mem[14530] = 198;
razn_h_mem[14531] = 74;
razn_h_mem[14532] = 204;
razn_h_mem[14533] = 80;
razn_h_mem[14534] = 210;
razn_h_mem[14535] = 86;
razn_h_mem[14536] = 216;
razn_h_mem[14537] = 92;
razn_h_mem[14538] = 222;
razn_h_mem[14539] = 98;
razn_h_mem[14540] = 228;
razn_h_mem[14541] = 104;
razn_h_mem[14542] = 234;
razn_h_mem[14543] = 110;
razn_h_mem[14544] = 240;
razn_h_mem[14545] = 116;
razn_h_mem[14546] = 246;
razn_h_mem[14547] = 122;
razn_h_mem[14548] = 252;
razn_h_mem[14549] = 128;
razn_h_mem[14550] = 4;
razn_h_mem[14551] = 134;
razn_h_mem[14552] = 10;
razn_h_mem[14553] = 140;
razn_h_mem[14554] = 16;
razn_h_mem[14555] = 146;
razn_h_mem[14556] = 22;
razn_h_mem[14557] = 152;
razn_h_mem[14558] = 28;
razn_h_mem[14559] = 158;
razn_h_mem[14560] = 34;
razn_h_mem[14561] = 164;
razn_h_mem[14562] = 40;
razn_h_mem[14563] = 170;
razn_h_mem[14564] = 46;
razn_h_mem[14565] = 176;
razn_h_mem[14566] = 52;
razn_h_mem[14567] = 182;
razn_h_mem[14568] = 58;
razn_h_mem[14569] = 188;
razn_h_mem[14570] = 64;
razn_h_mem[14571] = 194;
razn_h_mem[14572] = 70;
razn_h_mem[14573] = 200;
razn_h_mem[14574] = 76;
razn_h_mem[14575] = 206;
razn_h_mem[14576] = 82;
razn_h_mem[14577] = 212;
razn_h_mem[14578] = 88;
razn_h_mem[14579] = 218;
razn_h_mem[14580] = 94;
razn_h_mem[14581] = 224;
razn_h_mem[14582] = 100;
razn_h_mem[14583] = 230;
razn_h_mem[14584] = 106;
razn_h_mem[14585] = 236;
razn_h_mem[14586] = 112;
razn_h_mem[14587] = 242;
razn_h_mem[14588] = 118;
razn_h_mem[14589] = 248;
razn_h_mem[14590] = 124;
razn_h_mem[14591] = 255;
razn_h_mem[14592] = 0;
razn_h_mem[14593] = 130;
razn_h_mem[14594] = 6;
razn_h_mem[14595] = 136;
razn_h_mem[14596] = 12;
razn_h_mem[14597] = 142;
razn_h_mem[14598] = 18;
razn_h_mem[14599] = 148;
razn_h_mem[14600] = 24;
razn_h_mem[14601] = 154;
razn_h_mem[14602] = 30;
razn_h_mem[14603] = 160;
razn_h_mem[14604] = 36;
razn_h_mem[14605] = 166;
razn_h_mem[14606] = 42;
razn_h_mem[14607] = 172;
razn_h_mem[14608] = 48;
razn_h_mem[14609] = 178;
razn_h_mem[14610] = 54;
razn_h_mem[14611] = 184;
razn_h_mem[14612] = 60;
razn_h_mem[14613] = 190;
razn_h_mem[14614] = 66;
razn_h_mem[14615] = 196;
razn_h_mem[14616] = 72;
razn_h_mem[14617] = 202;
razn_h_mem[14618] = 78;
razn_h_mem[14619] = 208;
razn_h_mem[14620] = 84;
razn_h_mem[14621] = 214;
razn_h_mem[14622] = 90;
razn_h_mem[14623] = 220;
razn_h_mem[14624] = 96;
razn_h_mem[14625] = 226;
razn_h_mem[14626] = 102;
razn_h_mem[14627] = 232;
razn_h_mem[14628] = 108;
razn_h_mem[14629] = 238;
razn_h_mem[14630] = 114;
razn_h_mem[14631] = 244;
razn_h_mem[14632] = 120;
razn_h_mem[14633] = 250;
razn_h_mem[14634] = 126;
razn_h_mem[14635] = 2;
razn_h_mem[14636] = 132;
razn_h_mem[14637] = 8;
razn_h_mem[14638] = 138;
razn_h_mem[14639] = 14;
razn_h_mem[14640] = 144;
razn_h_mem[14641] = 20;
razn_h_mem[14642] = 150;
razn_h_mem[14643] = 26;
razn_h_mem[14644] = 156;
razn_h_mem[14645] = 32;
razn_h_mem[14646] = 162;
razn_h_mem[14647] = 38;
razn_h_mem[14648] = 168;
razn_h_mem[14649] = 44;
razn_h_mem[14650] = 174;
razn_h_mem[14651] = 50;
razn_h_mem[14652] = 180;
razn_h_mem[14653] = 56;
razn_h_mem[14654] = 186;
razn_h_mem[14655] = 62;
razn_h_mem[14656] = 192;
razn_h_mem[14657] = 68;
razn_h_mem[14658] = 198;
razn_h_mem[14659] = 74;
razn_h_mem[14660] = 204;
razn_h_mem[14661] = 80;
razn_h_mem[14662] = 210;
razn_h_mem[14663] = 86;
razn_h_mem[14664] = 216;
razn_h_mem[14665] = 92;
razn_h_mem[14666] = 222;
razn_h_mem[14667] = 98;
razn_h_mem[14668] = 228;
razn_h_mem[14669] = 104;
razn_h_mem[14670] = 234;
razn_h_mem[14671] = 110;
razn_h_mem[14672] = 240;
razn_h_mem[14673] = 116;
razn_h_mem[14674] = 246;
razn_h_mem[14675] = 122;
razn_h_mem[14676] = 252;
razn_h_mem[14677] = 128;
razn_h_mem[14678] = 4;
razn_h_mem[14679] = 134;
razn_h_mem[14680] = 10;
razn_h_mem[14681] = 140;
razn_h_mem[14682] = 16;
razn_h_mem[14683] = 146;
razn_h_mem[14684] = 22;
razn_h_mem[14685] = 152;
razn_h_mem[14686] = 28;
razn_h_mem[14687] = 158;
razn_h_mem[14688] = 34;
razn_h_mem[14689] = 164;
razn_h_mem[14690] = 40;
razn_h_mem[14691] = 170;
razn_h_mem[14692] = 46;
razn_h_mem[14693] = 176;
razn_h_mem[14694] = 52;
razn_h_mem[14695] = 182;
razn_h_mem[14696] = 58;
razn_h_mem[14697] = 188;
razn_h_mem[14698] = 64;
razn_h_mem[14699] = 194;
razn_h_mem[14700] = 70;
razn_h_mem[14701] = 200;
razn_h_mem[14702] = 76;
razn_h_mem[14703] = 206;
razn_h_mem[14704] = 82;
razn_h_mem[14705] = 212;
razn_h_mem[14706] = 88;
razn_h_mem[14707] = 218;
razn_h_mem[14708] = 94;
razn_h_mem[14709] = 224;
razn_h_mem[14710] = 100;
razn_h_mem[14711] = 230;
razn_h_mem[14712] = 106;
razn_h_mem[14713] = 236;
razn_h_mem[14714] = 112;
razn_h_mem[14715] = 242;
razn_h_mem[14716] = 118;
razn_h_mem[14717] = 248;
razn_h_mem[14718] = 124;
razn_h_mem[14719] = 255;
razn_h_mem[14720] = 0;
razn_h_mem[14721] = 130;
razn_h_mem[14722] = 6;
razn_h_mem[14723] = 136;
razn_h_mem[14724] = 12;
razn_h_mem[14725] = 142;
razn_h_mem[14726] = 18;
razn_h_mem[14727] = 148;
razn_h_mem[14728] = 24;
razn_h_mem[14729] = 154;
razn_h_mem[14730] = 30;
razn_h_mem[14731] = 160;
razn_h_mem[14732] = 36;
razn_h_mem[14733] = 166;
razn_h_mem[14734] = 42;
razn_h_mem[14735] = 172;
razn_h_mem[14736] = 48;
razn_h_mem[14737] = 178;
razn_h_mem[14738] = 54;
razn_h_mem[14739] = 184;
razn_h_mem[14740] = 60;
razn_h_mem[14741] = 190;
razn_h_mem[14742] = 66;
razn_h_mem[14743] = 196;
razn_h_mem[14744] = 72;
razn_h_mem[14745] = 202;
razn_h_mem[14746] = 78;
razn_h_mem[14747] = 208;
razn_h_mem[14748] = 84;
razn_h_mem[14749] = 214;
razn_h_mem[14750] = 90;
razn_h_mem[14751] = 220;
razn_h_mem[14752] = 96;
razn_h_mem[14753] = 226;
razn_h_mem[14754] = 102;
razn_h_mem[14755] = 232;
razn_h_mem[14756] = 108;
razn_h_mem[14757] = 238;
razn_h_mem[14758] = 114;
razn_h_mem[14759] = 244;
razn_h_mem[14760] = 120;
razn_h_mem[14761] = 250;
razn_h_mem[14762] = 126;
razn_h_mem[14763] = 2;
razn_h_mem[14764] = 132;
razn_h_mem[14765] = 8;
razn_h_mem[14766] = 138;
razn_h_mem[14767] = 14;
razn_h_mem[14768] = 144;
razn_h_mem[14769] = 20;
razn_h_mem[14770] = 150;
razn_h_mem[14771] = 26;
razn_h_mem[14772] = 156;
razn_h_mem[14773] = 32;
razn_h_mem[14774] = 162;
razn_h_mem[14775] = 38;
razn_h_mem[14776] = 168;
razn_h_mem[14777] = 44;
razn_h_mem[14778] = 174;
razn_h_mem[14779] = 50;
razn_h_mem[14780] = 180;
razn_h_mem[14781] = 56;
razn_h_mem[14782] = 186;
razn_h_mem[14783] = 62;
razn_h_mem[14784] = 192;
razn_h_mem[14785] = 68;
razn_h_mem[14786] = 198;
razn_h_mem[14787] = 74;
razn_h_mem[14788] = 204;
razn_h_mem[14789] = 80;
razn_h_mem[14790] = 210;
razn_h_mem[14791] = 86;
razn_h_mem[14792] = 216;
razn_h_mem[14793] = 92;
razn_h_mem[14794] = 222;
razn_h_mem[14795] = 98;
razn_h_mem[14796] = 228;
razn_h_mem[14797] = 104;
razn_h_mem[14798] = 234;
razn_h_mem[14799] = 110;
razn_h_mem[14800] = 240;
razn_h_mem[14801] = 116;
razn_h_mem[14802] = 246;
razn_h_mem[14803] = 122;
razn_h_mem[14804] = 252;
razn_h_mem[14805] = 128;
razn_h_mem[14806] = 4;
razn_h_mem[14807] = 134;
razn_h_mem[14808] = 10;
razn_h_mem[14809] = 140;
razn_h_mem[14810] = 16;
razn_h_mem[14811] = 146;
razn_h_mem[14812] = 22;
razn_h_mem[14813] = 152;
razn_h_mem[14814] = 28;
razn_h_mem[14815] = 158;
razn_h_mem[14816] = 34;
razn_h_mem[14817] = 164;
razn_h_mem[14818] = 40;
razn_h_mem[14819] = 170;
razn_h_mem[14820] = 46;
razn_h_mem[14821] = 176;
razn_h_mem[14822] = 52;
razn_h_mem[14823] = 182;
razn_h_mem[14824] = 58;
razn_h_mem[14825] = 188;
razn_h_mem[14826] = 64;
razn_h_mem[14827] = 194;
razn_h_mem[14828] = 70;
razn_h_mem[14829] = 200;
razn_h_mem[14830] = 76;
razn_h_mem[14831] = 206;
razn_h_mem[14832] = 82;
razn_h_mem[14833] = 212;
razn_h_mem[14834] = 88;
razn_h_mem[14835] = 218;
razn_h_mem[14836] = 94;
razn_h_mem[14837] = 224;
razn_h_mem[14838] = 100;
razn_h_mem[14839] = 230;
razn_h_mem[14840] = 106;
razn_h_mem[14841] = 236;
razn_h_mem[14842] = 112;
razn_h_mem[14843] = 242;
razn_h_mem[14844] = 118;
razn_h_mem[14845] = 248;
razn_h_mem[14846] = 124;
razn_h_mem[14847] = 255;
razn_h_mem[14848] = 0;
razn_h_mem[14849] = 130;
razn_h_mem[14850] = 6;
razn_h_mem[14851] = 136;
razn_h_mem[14852] = 12;
razn_h_mem[14853] = 142;
razn_h_mem[14854] = 18;
razn_h_mem[14855] = 148;
razn_h_mem[14856] = 24;
razn_h_mem[14857] = 154;
razn_h_mem[14858] = 30;
razn_h_mem[14859] = 160;
razn_h_mem[14860] = 36;
razn_h_mem[14861] = 166;
razn_h_mem[14862] = 42;
razn_h_mem[14863] = 172;
razn_h_mem[14864] = 48;
razn_h_mem[14865] = 178;
razn_h_mem[14866] = 54;
razn_h_mem[14867] = 184;
razn_h_mem[14868] = 60;
razn_h_mem[14869] = 190;
razn_h_mem[14870] = 66;
razn_h_mem[14871] = 196;
razn_h_mem[14872] = 72;
razn_h_mem[14873] = 202;
razn_h_mem[14874] = 78;
razn_h_mem[14875] = 208;
razn_h_mem[14876] = 84;
razn_h_mem[14877] = 214;
razn_h_mem[14878] = 90;
razn_h_mem[14879] = 220;
razn_h_mem[14880] = 96;
razn_h_mem[14881] = 226;
razn_h_mem[14882] = 102;
razn_h_mem[14883] = 232;
razn_h_mem[14884] = 108;
razn_h_mem[14885] = 238;
razn_h_mem[14886] = 114;
razn_h_mem[14887] = 244;
razn_h_mem[14888] = 120;
razn_h_mem[14889] = 250;
razn_h_mem[14890] = 126;
razn_h_mem[14891] = 2;
razn_h_mem[14892] = 132;
razn_h_mem[14893] = 8;
razn_h_mem[14894] = 138;
razn_h_mem[14895] = 14;
razn_h_mem[14896] = 144;
razn_h_mem[14897] = 20;
razn_h_mem[14898] = 150;
razn_h_mem[14899] = 26;
razn_h_mem[14900] = 156;
razn_h_mem[14901] = 32;
razn_h_mem[14902] = 162;
razn_h_mem[14903] = 38;
razn_h_mem[14904] = 168;
razn_h_mem[14905] = 44;
razn_h_mem[14906] = 174;
razn_h_mem[14907] = 50;
razn_h_mem[14908] = 180;
razn_h_mem[14909] = 56;
razn_h_mem[14910] = 186;
razn_h_mem[14911] = 62;
razn_h_mem[14912] = 192;
razn_h_mem[14913] = 68;
razn_h_mem[14914] = 198;
razn_h_mem[14915] = 74;
razn_h_mem[14916] = 204;
razn_h_mem[14917] = 80;
razn_h_mem[14918] = 210;
razn_h_mem[14919] = 86;
razn_h_mem[14920] = 216;
razn_h_mem[14921] = 92;
razn_h_mem[14922] = 222;
razn_h_mem[14923] = 98;
razn_h_mem[14924] = 228;
razn_h_mem[14925] = 104;
razn_h_mem[14926] = 234;
razn_h_mem[14927] = 110;
razn_h_mem[14928] = 240;
razn_h_mem[14929] = 116;
razn_h_mem[14930] = 246;
razn_h_mem[14931] = 122;
razn_h_mem[14932] = 252;
razn_h_mem[14933] = 128;
razn_h_mem[14934] = 4;
razn_h_mem[14935] = 134;
razn_h_mem[14936] = 10;
razn_h_mem[14937] = 140;
razn_h_mem[14938] = 16;
razn_h_mem[14939] = 146;
razn_h_mem[14940] = 22;
razn_h_mem[14941] = 152;
razn_h_mem[14942] = 28;
razn_h_mem[14943] = 158;
razn_h_mem[14944] = 34;
razn_h_mem[14945] = 164;
razn_h_mem[14946] = 40;
razn_h_mem[14947] = 170;
razn_h_mem[14948] = 46;
razn_h_mem[14949] = 176;
razn_h_mem[14950] = 52;
razn_h_mem[14951] = 182;
razn_h_mem[14952] = 58;
razn_h_mem[14953] = 188;
razn_h_mem[14954] = 64;
razn_h_mem[14955] = 194;
razn_h_mem[14956] = 70;
razn_h_mem[14957] = 200;
razn_h_mem[14958] = 76;
razn_h_mem[14959] = 206;
razn_h_mem[14960] = 82;
razn_h_mem[14961] = 212;
razn_h_mem[14962] = 88;
razn_h_mem[14963] = 218;
razn_h_mem[14964] = 94;
razn_h_mem[14965] = 224;
razn_h_mem[14966] = 100;
razn_h_mem[14967] = 230;
razn_h_mem[14968] = 106;
razn_h_mem[14969] = 236;
razn_h_mem[14970] = 112;
razn_h_mem[14971] = 242;
razn_h_mem[14972] = 118;
razn_h_mem[14973] = 248;
razn_h_mem[14974] = 124;
razn_h_mem[14975] = 255;
razn_h_mem[14976] = 0;
razn_h_mem[14977] = 130;
razn_h_mem[14978] = 6;
razn_h_mem[14979] = 136;
razn_h_mem[14980] = 12;
razn_h_mem[14981] = 142;
razn_h_mem[14982] = 18;
razn_h_mem[14983] = 148;
razn_h_mem[14984] = 24;
razn_h_mem[14985] = 154;
razn_h_mem[14986] = 30;
razn_h_mem[14987] = 160;
razn_h_mem[14988] = 36;
razn_h_mem[14989] = 166;
razn_h_mem[14990] = 42;
razn_h_mem[14991] = 172;
razn_h_mem[14992] = 48;
razn_h_mem[14993] = 178;
razn_h_mem[14994] = 54;
razn_h_mem[14995] = 184;
razn_h_mem[14996] = 60;
razn_h_mem[14997] = 190;
razn_h_mem[14998] = 66;
razn_h_mem[14999] = 196;
razn_h_mem[15000] = 72;
razn_h_mem[15001] = 202;
razn_h_mem[15002] = 78;
razn_h_mem[15003] = 208;
razn_h_mem[15004] = 84;
razn_h_mem[15005] = 214;
razn_h_mem[15006] = 90;
razn_h_mem[15007] = 220;
razn_h_mem[15008] = 96;
razn_h_mem[15009] = 226;
razn_h_mem[15010] = 102;
razn_h_mem[15011] = 232;
razn_h_mem[15012] = 108;
razn_h_mem[15013] = 238;
razn_h_mem[15014] = 114;
razn_h_mem[15015] = 244;
razn_h_mem[15016] = 120;
razn_h_mem[15017] = 250;
razn_h_mem[15018] = 126;
razn_h_mem[15019] = 2;
razn_h_mem[15020] = 132;
razn_h_mem[15021] = 8;
razn_h_mem[15022] = 138;
razn_h_mem[15023] = 14;
razn_h_mem[15024] = 144;
razn_h_mem[15025] = 20;
razn_h_mem[15026] = 150;
razn_h_mem[15027] = 26;
razn_h_mem[15028] = 156;
razn_h_mem[15029] = 32;
razn_h_mem[15030] = 162;
razn_h_mem[15031] = 38;
razn_h_mem[15032] = 168;
razn_h_mem[15033] = 44;
razn_h_mem[15034] = 174;
razn_h_mem[15035] = 50;
razn_h_mem[15036] = 180;
razn_h_mem[15037] = 56;
razn_h_mem[15038] = 186;
razn_h_mem[15039] = 62;
razn_h_mem[15040] = 192;
razn_h_mem[15041] = 68;
razn_h_mem[15042] = 198;
razn_h_mem[15043] = 74;
razn_h_mem[15044] = 204;
razn_h_mem[15045] = 80;
razn_h_mem[15046] = 210;
razn_h_mem[15047] = 86;
razn_h_mem[15048] = 216;
razn_h_mem[15049] = 92;
razn_h_mem[15050] = 222;
razn_h_mem[15051] = 98;
razn_h_mem[15052] = 228;
razn_h_mem[15053] = 104;
razn_h_mem[15054] = 234;
razn_h_mem[15055] = 110;
razn_h_mem[15056] = 240;
razn_h_mem[15057] = 116;
razn_h_mem[15058] = 246;
razn_h_mem[15059] = 122;
razn_h_mem[15060] = 252;
razn_h_mem[15061] = 128;
razn_h_mem[15062] = 4;
razn_h_mem[15063] = 134;
razn_h_mem[15064] = 10;
razn_h_mem[15065] = 140;
razn_h_mem[15066] = 16;
razn_h_mem[15067] = 146;
razn_h_mem[15068] = 22;
razn_h_mem[15069] = 152;
razn_h_mem[15070] = 28;
razn_h_mem[15071] = 158;
razn_h_mem[15072] = 34;
razn_h_mem[15073] = 164;
razn_h_mem[15074] = 40;
razn_h_mem[15075] = 170;
razn_h_mem[15076] = 46;
razn_h_mem[15077] = 176;
razn_h_mem[15078] = 52;
razn_h_mem[15079] = 182;
razn_h_mem[15080] = 58;
razn_h_mem[15081] = 188;
razn_h_mem[15082] = 64;
razn_h_mem[15083] = 194;
razn_h_mem[15084] = 70;
razn_h_mem[15085] = 200;
razn_h_mem[15086] = 76;
razn_h_mem[15087] = 206;
razn_h_mem[15088] = 82;
razn_h_mem[15089] = 212;
razn_h_mem[15090] = 88;
razn_h_mem[15091] = 218;
razn_h_mem[15092] = 94;
razn_h_mem[15093] = 224;
razn_h_mem[15094] = 100;
razn_h_mem[15095] = 230;
razn_h_mem[15096] = 106;
razn_h_mem[15097] = 236;
razn_h_mem[15098] = 112;
razn_h_mem[15099] = 242;
razn_h_mem[15100] = 118;
razn_h_mem[15101] = 248;
razn_h_mem[15102] = 124;
razn_h_mem[15103] = 255;
razn_h_mem[15104] = 0;
razn_h_mem[15105] = 130;
razn_h_mem[15106] = 6;
razn_h_mem[15107] = 136;
razn_h_mem[15108] = 12;
razn_h_mem[15109] = 142;
razn_h_mem[15110] = 18;
razn_h_mem[15111] = 148;
razn_h_mem[15112] = 24;
razn_h_mem[15113] = 154;
razn_h_mem[15114] = 30;
razn_h_mem[15115] = 160;
razn_h_mem[15116] = 36;
razn_h_mem[15117] = 166;
razn_h_mem[15118] = 42;
razn_h_mem[15119] = 172;
razn_h_mem[15120] = 48;
razn_h_mem[15121] = 178;
razn_h_mem[15122] = 54;
razn_h_mem[15123] = 184;
razn_h_mem[15124] = 60;
razn_h_mem[15125] = 190;
razn_h_mem[15126] = 66;
razn_h_mem[15127] = 196;
razn_h_mem[15128] = 72;
razn_h_mem[15129] = 202;
razn_h_mem[15130] = 78;
razn_h_mem[15131] = 208;
razn_h_mem[15132] = 84;
razn_h_mem[15133] = 214;
razn_h_mem[15134] = 90;
razn_h_mem[15135] = 220;
razn_h_mem[15136] = 96;
razn_h_mem[15137] = 226;
razn_h_mem[15138] = 102;
razn_h_mem[15139] = 232;
razn_h_mem[15140] = 108;
razn_h_mem[15141] = 238;
razn_h_mem[15142] = 114;
razn_h_mem[15143] = 244;
razn_h_mem[15144] = 120;
razn_h_mem[15145] = 250;
razn_h_mem[15146] = 126;
razn_h_mem[15147] = 2;
razn_h_mem[15148] = 132;
razn_h_mem[15149] = 8;
razn_h_mem[15150] = 138;
razn_h_mem[15151] = 14;
razn_h_mem[15152] = 144;
razn_h_mem[15153] = 20;
razn_h_mem[15154] = 150;
razn_h_mem[15155] = 26;
razn_h_mem[15156] = 156;
razn_h_mem[15157] = 32;
razn_h_mem[15158] = 162;
razn_h_mem[15159] = 38;
razn_h_mem[15160] = 168;
razn_h_mem[15161] = 44;
razn_h_mem[15162] = 174;
razn_h_mem[15163] = 50;
razn_h_mem[15164] = 180;
razn_h_mem[15165] = 56;
razn_h_mem[15166] = 186;
razn_h_mem[15167] = 62;
razn_h_mem[15168] = 192;
razn_h_mem[15169] = 68;
razn_h_mem[15170] = 198;
razn_h_mem[15171] = 74;
razn_h_mem[15172] = 204;
razn_h_mem[15173] = 80;
razn_h_mem[15174] = 210;
razn_h_mem[15175] = 86;
razn_h_mem[15176] = 216;
razn_h_mem[15177] = 92;
razn_h_mem[15178] = 222;
razn_h_mem[15179] = 98;
razn_h_mem[15180] = 228;
razn_h_mem[15181] = 104;
razn_h_mem[15182] = 234;
razn_h_mem[15183] = 110;
razn_h_mem[15184] = 240;
razn_h_mem[15185] = 116;
razn_h_mem[15186] = 246;
razn_h_mem[15187] = 122;
razn_h_mem[15188] = 252;
razn_h_mem[15189] = 128;
razn_h_mem[15190] = 4;
razn_h_mem[15191] = 134;
razn_h_mem[15192] = 10;
razn_h_mem[15193] = 140;
razn_h_mem[15194] = 16;
razn_h_mem[15195] = 146;
razn_h_mem[15196] = 22;
razn_h_mem[15197] = 152;
razn_h_mem[15198] = 28;
razn_h_mem[15199] = 158;
razn_h_mem[15200] = 34;
razn_h_mem[15201] = 164;
razn_h_mem[15202] = 40;
razn_h_mem[15203] = 170;
razn_h_mem[15204] = 46;
razn_h_mem[15205] = 176;
razn_h_mem[15206] = 52;
razn_h_mem[15207] = 182;
razn_h_mem[15208] = 58;
razn_h_mem[15209] = 188;
razn_h_mem[15210] = 64;
razn_h_mem[15211] = 194;
razn_h_mem[15212] = 70;
razn_h_mem[15213] = 200;
razn_h_mem[15214] = 76;
razn_h_mem[15215] = 206;
razn_h_mem[15216] = 82;
razn_h_mem[15217] = 212;
razn_h_mem[15218] = 88;
razn_h_mem[15219] = 218;
razn_h_mem[15220] = 94;
razn_h_mem[15221] = 224;
razn_h_mem[15222] = 100;
razn_h_mem[15223] = 230;
razn_h_mem[15224] = 106;
razn_h_mem[15225] = 236;
razn_h_mem[15226] = 112;
razn_h_mem[15227] = 242;
razn_h_mem[15228] = 118;
razn_h_mem[15229] = 248;
razn_h_mem[15230] = 124;
razn_h_mem[15231] = 255;
razn_h_mem[15232] = 0;
razn_h_mem[15233] = 130;
razn_h_mem[15234] = 6;
razn_h_mem[15235] = 136;
razn_h_mem[15236] = 12;
razn_h_mem[15237] = 142;
razn_h_mem[15238] = 18;
razn_h_mem[15239] = 148;
razn_h_mem[15240] = 24;
razn_h_mem[15241] = 154;
razn_h_mem[15242] = 30;
razn_h_mem[15243] = 160;
razn_h_mem[15244] = 36;
razn_h_mem[15245] = 166;
razn_h_mem[15246] = 42;
razn_h_mem[15247] = 172;
razn_h_mem[15248] = 48;
razn_h_mem[15249] = 178;
razn_h_mem[15250] = 54;
razn_h_mem[15251] = 184;
razn_h_mem[15252] = 60;
razn_h_mem[15253] = 190;
razn_h_mem[15254] = 66;
razn_h_mem[15255] = 196;
razn_h_mem[15256] = 72;
razn_h_mem[15257] = 202;
razn_h_mem[15258] = 78;
razn_h_mem[15259] = 208;
razn_h_mem[15260] = 84;
razn_h_mem[15261] = 214;
razn_h_mem[15262] = 90;
razn_h_mem[15263] = 220;
razn_h_mem[15264] = 96;
razn_h_mem[15265] = 226;
razn_h_mem[15266] = 102;
razn_h_mem[15267] = 232;
razn_h_mem[15268] = 108;
razn_h_mem[15269] = 238;
razn_h_mem[15270] = 114;
razn_h_mem[15271] = 244;
razn_h_mem[15272] = 120;
razn_h_mem[15273] = 250;
razn_h_mem[15274] = 126;
razn_h_mem[15275] = 2;
razn_h_mem[15276] = 132;
razn_h_mem[15277] = 8;
razn_h_mem[15278] = 138;
razn_h_mem[15279] = 14;
razn_h_mem[15280] = 144;
razn_h_mem[15281] = 20;
razn_h_mem[15282] = 150;
razn_h_mem[15283] = 26;
razn_h_mem[15284] = 156;
razn_h_mem[15285] = 32;
razn_h_mem[15286] = 162;
razn_h_mem[15287] = 38;
razn_h_mem[15288] = 168;
razn_h_mem[15289] = 44;
razn_h_mem[15290] = 174;
razn_h_mem[15291] = 50;
razn_h_mem[15292] = 180;
razn_h_mem[15293] = 56;
razn_h_mem[15294] = 186;
razn_h_mem[15295] = 62;
razn_h_mem[15296] = 192;
razn_h_mem[15297] = 68;
razn_h_mem[15298] = 198;
razn_h_mem[15299] = 74;
razn_h_mem[15300] = 204;
razn_h_mem[15301] = 80;
razn_h_mem[15302] = 210;
razn_h_mem[15303] = 86;
razn_h_mem[15304] = 216;
razn_h_mem[15305] = 92;
razn_h_mem[15306] = 222;
razn_h_mem[15307] = 98;
razn_h_mem[15308] = 228;
razn_h_mem[15309] = 104;
razn_h_mem[15310] = 234;
razn_h_mem[15311] = 110;
razn_h_mem[15312] = 240;
razn_h_mem[15313] = 116;
razn_h_mem[15314] = 246;
razn_h_mem[15315] = 122;
razn_h_mem[15316] = 252;
razn_h_mem[15317] = 128;
razn_h_mem[15318] = 4;
razn_h_mem[15319] = 134;
razn_h_mem[15320] = 10;
razn_h_mem[15321] = 140;
razn_h_mem[15322] = 16;
razn_h_mem[15323] = 146;
razn_h_mem[15324] = 22;
razn_h_mem[15325] = 152;
razn_h_mem[15326] = 28;
razn_h_mem[15327] = 158;
razn_h_mem[15328] = 34;
razn_h_mem[15329] = 164;
razn_h_mem[15330] = 40;
razn_h_mem[15331] = 170;
razn_h_mem[15332] = 46;
razn_h_mem[15333] = 176;
razn_h_mem[15334] = 52;
razn_h_mem[15335] = 182;
razn_h_mem[15336] = 58;
razn_h_mem[15337] = 188;
razn_h_mem[15338] = 64;
razn_h_mem[15339] = 194;
razn_h_mem[15340] = 70;
razn_h_mem[15341] = 200;
razn_h_mem[15342] = 76;
razn_h_mem[15343] = 206;
razn_h_mem[15344] = 82;
razn_h_mem[15345] = 212;
razn_h_mem[15346] = 88;
razn_h_mem[15347] = 218;
razn_h_mem[15348] = 94;
razn_h_mem[15349] = 224;
razn_h_mem[15350] = 100;
razn_h_mem[15351] = 230;
razn_h_mem[15352] = 106;
razn_h_mem[15353] = 236;
razn_h_mem[15354] = 112;
razn_h_mem[15355] = 242;
razn_h_mem[15356] = 118;
razn_h_mem[15357] = 248;
razn_h_mem[15358] = 124;
razn_h_mem[15359] = 255;
razn_h_mem[15360] = 0;
razn_h_mem[15361] = 130;
razn_h_mem[15362] = 6;
razn_h_mem[15363] = 136;
razn_h_mem[15364] = 12;
razn_h_mem[15365] = 142;
razn_h_mem[15366] = 18;
razn_h_mem[15367] = 148;
razn_h_mem[15368] = 24;
razn_h_mem[15369] = 154;
razn_h_mem[15370] = 30;
razn_h_mem[15371] = 160;
razn_h_mem[15372] = 36;
razn_h_mem[15373] = 166;
razn_h_mem[15374] = 42;
razn_h_mem[15375] = 172;
razn_h_mem[15376] = 48;
razn_h_mem[15377] = 178;
razn_h_mem[15378] = 54;
razn_h_mem[15379] = 184;
razn_h_mem[15380] = 60;
razn_h_mem[15381] = 190;
razn_h_mem[15382] = 66;
razn_h_mem[15383] = 196;
razn_h_mem[15384] = 72;
razn_h_mem[15385] = 202;
razn_h_mem[15386] = 78;
razn_h_mem[15387] = 208;
razn_h_mem[15388] = 84;
razn_h_mem[15389] = 214;
razn_h_mem[15390] = 90;
razn_h_mem[15391] = 220;
razn_h_mem[15392] = 96;
razn_h_mem[15393] = 226;
razn_h_mem[15394] = 102;
razn_h_mem[15395] = 232;
razn_h_mem[15396] = 108;
razn_h_mem[15397] = 238;
razn_h_mem[15398] = 114;
razn_h_mem[15399] = 244;
razn_h_mem[15400] = 120;
razn_h_mem[15401] = 250;
razn_h_mem[15402] = 126;
razn_h_mem[15403] = 2;
razn_h_mem[15404] = 132;
razn_h_mem[15405] = 8;
razn_h_mem[15406] = 138;
razn_h_mem[15407] = 14;
razn_h_mem[15408] = 144;
razn_h_mem[15409] = 20;
razn_h_mem[15410] = 150;
razn_h_mem[15411] = 26;
razn_h_mem[15412] = 156;
razn_h_mem[15413] = 32;
razn_h_mem[15414] = 162;
razn_h_mem[15415] = 38;
razn_h_mem[15416] = 168;
razn_h_mem[15417] = 44;
razn_h_mem[15418] = 174;
razn_h_mem[15419] = 50;
razn_h_mem[15420] = 180;
razn_h_mem[15421] = 56;
razn_h_mem[15422] = 186;
razn_h_mem[15423] = 62;
razn_h_mem[15424] = 192;
razn_h_mem[15425] = 68;
razn_h_mem[15426] = 198;
razn_h_mem[15427] = 74;
razn_h_mem[15428] = 204;
razn_h_mem[15429] = 80;
razn_h_mem[15430] = 210;
razn_h_mem[15431] = 86;
razn_h_mem[15432] = 216;
razn_h_mem[15433] = 92;
razn_h_mem[15434] = 222;
razn_h_mem[15435] = 98;
razn_h_mem[15436] = 228;
razn_h_mem[15437] = 104;
razn_h_mem[15438] = 234;
razn_h_mem[15439] = 110;
razn_h_mem[15440] = 240;
razn_h_mem[15441] = 116;
razn_h_mem[15442] = 246;
razn_h_mem[15443] = 122;
razn_h_mem[15444] = 252;
razn_h_mem[15445] = 128;
razn_h_mem[15446] = 4;
razn_h_mem[15447] = 134;
razn_h_mem[15448] = 10;
razn_h_mem[15449] = 140;
razn_h_mem[15450] = 16;
razn_h_mem[15451] = 146;
razn_h_mem[15452] = 22;
razn_h_mem[15453] = 152;
razn_h_mem[15454] = 28;
razn_h_mem[15455] = 158;
razn_h_mem[15456] = 34;
razn_h_mem[15457] = 164;
razn_h_mem[15458] = 40;
razn_h_mem[15459] = 170;
razn_h_mem[15460] = 46;
razn_h_mem[15461] = 176;
razn_h_mem[15462] = 52;
razn_h_mem[15463] = 182;
razn_h_mem[15464] = 58;
razn_h_mem[15465] = 188;
razn_h_mem[15466] = 64;
razn_h_mem[15467] = 194;
razn_h_mem[15468] = 70;
razn_h_mem[15469] = 200;
razn_h_mem[15470] = 76;
razn_h_mem[15471] = 206;
razn_h_mem[15472] = 82;
razn_h_mem[15473] = 212;
razn_h_mem[15474] = 88;
razn_h_mem[15475] = 218;
razn_h_mem[15476] = 94;
razn_h_mem[15477] = 224;
razn_h_mem[15478] = 100;
razn_h_mem[15479] = 230;
razn_h_mem[15480] = 106;
razn_h_mem[15481] = 236;
razn_h_mem[15482] = 112;
razn_h_mem[15483] = 242;
razn_h_mem[15484] = 118;
razn_h_mem[15485] = 248;
razn_h_mem[15486] = 124;
razn_h_mem[15487] = 255;
razn_h_mem[15488] = 0;
razn_h_mem[15489] = 130;
razn_h_mem[15490] = 6;
razn_h_mem[15491] = 136;
razn_h_mem[15492] = 12;
razn_h_mem[15493] = 142;
razn_h_mem[15494] = 18;
razn_h_mem[15495] = 148;
razn_h_mem[15496] = 24;
razn_h_mem[15497] = 154;
razn_h_mem[15498] = 30;
razn_h_mem[15499] = 160;
razn_h_mem[15500] = 36;
razn_h_mem[15501] = 166;
razn_h_mem[15502] = 42;
razn_h_mem[15503] = 172;
razn_h_mem[15504] = 48;
razn_h_mem[15505] = 178;
razn_h_mem[15506] = 54;
razn_h_mem[15507] = 184;
razn_h_mem[15508] = 60;
razn_h_mem[15509] = 190;
razn_h_mem[15510] = 66;
razn_h_mem[15511] = 196;
razn_h_mem[15512] = 72;
razn_h_mem[15513] = 202;
razn_h_mem[15514] = 78;
razn_h_mem[15515] = 208;
razn_h_mem[15516] = 84;
razn_h_mem[15517] = 214;
razn_h_mem[15518] = 90;
razn_h_mem[15519] = 220;
razn_h_mem[15520] = 96;
razn_h_mem[15521] = 226;
razn_h_mem[15522] = 102;
razn_h_mem[15523] = 232;
razn_h_mem[15524] = 108;
razn_h_mem[15525] = 238;
razn_h_mem[15526] = 114;
razn_h_mem[15527] = 244;
razn_h_mem[15528] = 120;
razn_h_mem[15529] = 250;
razn_h_mem[15530] = 126;
razn_h_mem[15531] = 2;
razn_h_mem[15532] = 132;
razn_h_mem[15533] = 8;
razn_h_mem[15534] = 138;
razn_h_mem[15535] = 14;
razn_h_mem[15536] = 144;
razn_h_mem[15537] = 20;
razn_h_mem[15538] = 150;
razn_h_mem[15539] = 26;
razn_h_mem[15540] = 156;
razn_h_mem[15541] = 32;
razn_h_mem[15542] = 162;
razn_h_mem[15543] = 38;
razn_h_mem[15544] = 168;
razn_h_mem[15545] = 44;
razn_h_mem[15546] = 174;
razn_h_mem[15547] = 50;
razn_h_mem[15548] = 180;
razn_h_mem[15549] = 56;
razn_h_mem[15550] = 186;
razn_h_mem[15551] = 62;
razn_h_mem[15552] = 192;
razn_h_mem[15553] = 68;
razn_h_mem[15554] = 198;
razn_h_mem[15555] = 74;
razn_h_mem[15556] = 204;
razn_h_mem[15557] = 80;
razn_h_mem[15558] = 210;
razn_h_mem[15559] = 86;
razn_h_mem[15560] = 216;
razn_h_mem[15561] = 92;
razn_h_mem[15562] = 222;
razn_h_mem[15563] = 98;
razn_h_mem[15564] = 228;
razn_h_mem[15565] = 104;
razn_h_mem[15566] = 234;
razn_h_mem[15567] = 110;
razn_h_mem[15568] = 240;
razn_h_mem[15569] = 116;
razn_h_mem[15570] = 246;
razn_h_mem[15571] = 122;
razn_h_mem[15572] = 252;
razn_h_mem[15573] = 128;
razn_h_mem[15574] = 4;
razn_h_mem[15575] = 134;
razn_h_mem[15576] = 10;
razn_h_mem[15577] = 140;
razn_h_mem[15578] = 16;
razn_h_mem[15579] = 146;
razn_h_mem[15580] = 22;
razn_h_mem[15581] = 152;
razn_h_mem[15582] = 28;
razn_h_mem[15583] = 158;
razn_h_mem[15584] = 34;
razn_h_mem[15585] = 164;
razn_h_mem[15586] = 40;
razn_h_mem[15587] = 170;
razn_h_mem[15588] = 46;
razn_h_mem[15589] = 176;
razn_h_mem[15590] = 52;
razn_h_mem[15591] = 182;
razn_h_mem[15592] = 58;
razn_h_mem[15593] = 188;
razn_h_mem[15594] = 64;
razn_h_mem[15595] = 194;
razn_h_mem[15596] = 70;
razn_h_mem[15597] = 200;
razn_h_mem[15598] = 76;
razn_h_mem[15599] = 206;
razn_h_mem[15600] = 82;
razn_h_mem[15601] = 212;
razn_h_mem[15602] = 88;
razn_h_mem[15603] = 218;
razn_h_mem[15604] = 94;
razn_h_mem[15605] = 224;
razn_h_mem[15606] = 100;
razn_h_mem[15607] = 230;
razn_h_mem[15608] = 106;
razn_h_mem[15609] = 236;
razn_h_mem[15610] = 112;
razn_h_mem[15611] = 242;
razn_h_mem[15612] = 118;
razn_h_mem[15613] = 248;
razn_h_mem[15614] = 124;
razn_h_mem[15615] = 255;
razn_h_mem[15616] = 0;
razn_h_mem[15617] = 130;
razn_h_mem[15618] = 6;
razn_h_mem[15619] = 136;
razn_h_mem[15620] = 12;
razn_h_mem[15621] = 142;
razn_h_mem[15622] = 18;
razn_h_mem[15623] = 148;
razn_h_mem[15624] = 24;
razn_h_mem[15625] = 154;
razn_h_mem[15626] = 30;
razn_h_mem[15627] = 160;
razn_h_mem[15628] = 36;
razn_h_mem[15629] = 166;
razn_h_mem[15630] = 42;
razn_h_mem[15631] = 172;
razn_h_mem[15632] = 48;
razn_h_mem[15633] = 178;
razn_h_mem[15634] = 54;
razn_h_mem[15635] = 184;
razn_h_mem[15636] = 60;
razn_h_mem[15637] = 190;
razn_h_mem[15638] = 66;
razn_h_mem[15639] = 196;
razn_h_mem[15640] = 72;
razn_h_mem[15641] = 202;
razn_h_mem[15642] = 78;
razn_h_mem[15643] = 208;
razn_h_mem[15644] = 84;
razn_h_mem[15645] = 214;
razn_h_mem[15646] = 90;
razn_h_mem[15647] = 220;
razn_h_mem[15648] = 96;
razn_h_mem[15649] = 226;
razn_h_mem[15650] = 102;
razn_h_mem[15651] = 232;
razn_h_mem[15652] = 108;
razn_h_mem[15653] = 238;
razn_h_mem[15654] = 114;
razn_h_mem[15655] = 244;
razn_h_mem[15656] = 120;
razn_h_mem[15657] = 250;
razn_h_mem[15658] = 126;
razn_h_mem[15659] = 2;
razn_h_mem[15660] = 132;
razn_h_mem[15661] = 8;
razn_h_mem[15662] = 138;
razn_h_mem[15663] = 14;
razn_h_mem[15664] = 144;
razn_h_mem[15665] = 20;
razn_h_mem[15666] = 150;
razn_h_mem[15667] = 26;
razn_h_mem[15668] = 156;
razn_h_mem[15669] = 32;
razn_h_mem[15670] = 162;
razn_h_mem[15671] = 38;
razn_h_mem[15672] = 168;
razn_h_mem[15673] = 44;
razn_h_mem[15674] = 174;
razn_h_mem[15675] = 50;
razn_h_mem[15676] = 180;
razn_h_mem[15677] = 56;
razn_h_mem[15678] = 186;
razn_h_mem[15679] = 62;
razn_h_mem[15680] = 192;
razn_h_mem[15681] = 68;
razn_h_mem[15682] = 198;
razn_h_mem[15683] = 74;
razn_h_mem[15684] = 204;
razn_h_mem[15685] = 80;
razn_h_mem[15686] = 210;
razn_h_mem[15687] = 86;
razn_h_mem[15688] = 216;
razn_h_mem[15689] = 92;
razn_h_mem[15690] = 222;
razn_h_mem[15691] = 98;
razn_h_mem[15692] = 228;
razn_h_mem[15693] = 104;
razn_h_mem[15694] = 234;
razn_h_mem[15695] = 110;
razn_h_mem[15696] = 240;
razn_h_mem[15697] = 116;
razn_h_mem[15698] = 246;
razn_h_mem[15699] = 122;
razn_h_mem[15700] = 252;
razn_h_mem[15701] = 128;
razn_h_mem[15702] = 4;
razn_h_mem[15703] = 134;
razn_h_mem[15704] = 10;
razn_h_mem[15705] = 140;
razn_h_mem[15706] = 16;
razn_h_mem[15707] = 146;
razn_h_mem[15708] = 22;
razn_h_mem[15709] = 152;
razn_h_mem[15710] = 28;
razn_h_mem[15711] = 158;
razn_h_mem[15712] = 34;
razn_h_mem[15713] = 164;
razn_h_mem[15714] = 40;
razn_h_mem[15715] = 170;
razn_h_mem[15716] = 46;
razn_h_mem[15717] = 176;
razn_h_mem[15718] = 52;
razn_h_mem[15719] = 182;
razn_h_mem[15720] = 58;
razn_h_mem[15721] = 188;
razn_h_mem[15722] = 64;
razn_h_mem[15723] = 194;
razn_h_mem[15724] = 70;
razn_h_mem[15725] = 200;
razn_h_mem[15726] = 76;
razn_h_mem[15727] = 206;
razn_h_mem[15728] = 82;
razn_h_mem[15729] = 212;
razn_h_mem[15730] = 88;
razn_h_mem[15731] = 218;
razn_h_mem[15732] = 94;
razn_h_mem[15733] = 224;
razn_h_mem[15734] = 100;
razn_h_mem[15735] = 230;
razn_h_mem[15736] = 106;
razn_h_mem[15737] = 236;
razn_h_mem[15738] = 112;
razn_h_mem[15739] = 242;
razn_h_mem[15740] = 118;
razn_h_mem[15741] = 248;
razn_h_mem[15742] = 124;
razn_h_mem[15743] = 255;
razn_h_mem[15744] = 0;
razn_h_mem[15745] = 130;
razn_h_mem[15746] = 6;
razn_h_mem[15747] = 136;
razn_h_mem[15748] = 12;
razn_h_mem[15749] = 142;
razn_h_mem[15750] = 18;
razn_h_mem[15751] = 148;
razn_h_mem[15752] = 24;
razn_h_mem[15753] = 154;
razn_h_mem[15754] = 30;
razn_h_mem[15755] = 160;
razn_h_mem[15756] = 36;
razn_h_mem[15757] = 166;
razn_h_mem[15758] = 42;
razn_h_mem[15759] = 172;
razn_h_mem[15760] = 48;
razn_h_mem[15761] = 178;
razn_h_mem[15762] = 54;
razn_h_mem[15763] = 184;
razn_h_mem[15764] = 60;
razn_h_mem[15765] = 190;
razn_h_mem[15766] = 66;
razn_h_mem[15767] = 196;
razn_h_mem[15768] = 72;
razn_h_mem[15769] = 202;
razn_h_mem[15770] = 78;
razn_h_mem[15771] = 208;
razn_h_mem[15772] = 84;
razn_h_mem[15773] = 214;
razn_h_mem[15774] = 90;
razn_h_mem[15775] = 220;
razn_h_mem[15776] = 96;
razn_h_mem[15777] = 226;
razn_h_mem[15778] = 102;
razn_h_mem[15779] = 232;
razn_h_mem[15780] = 108;
razn_h_mem[15781] = 238;
razn_h_mem[15782] = 114;
razn_h_mem[15783] = 244;
razn_h_mem[15784] = 120;
razn_h_mem[15785] = 250;
razn_h_mem[15786] = 126;
razn_h_mem[15787] = 2;
razn_h_mem[15788] = 132;
razn_h_mem[15789] = 8;
razn_h_mem[15790] = 138;
razn_h_mem[15791] = 14;
razn_h_mem[15792] = 144;
razn_h_mem[15793] = 20;
razn_h_mem[15794] = 150;
razn_h_mem[15795] = 26;
razn_h_mem[15796] = 156;
razn_h_mem[15797] = 32;
razn_h_mem[15798] = 162;
razn_h_mem[15799] = 38;
razn_h_mem[15800] = 168;
razn_h_mem[15801] = 44;
razn_h_mem[15802] = 174;
razn_h_mem[15803] = 50;
razn_h_mem[15804] = 180;
razn_h_mem[15805] = 56;
razn_h_mem[15806] = 186;
razn_h_mem[15807] = 62;
razn_h_mem[15808] = 192;
razn_h_mem[15809] = 68;
razn_h_mem[15810] = 198;
razn_h_mem[15811] = 74;
razn_h_mem[15812] = 204;
razn_h_mem[15813] = 80;
razn_h_mem[15814] = 210;
razn_h_mem[15815] = 86;
razn_h_mem[15816] = 216;
razn_h_mem[15817] = 92;
razn_h_mem[15818] = 222;
razn_h_mem[15819] = 98;
razn_h_mem[15820] = 228;
razn_h_mem[15821] = 104;
razn_h_mem[15822] = 234;
razn_h_mem[15823] = 110;
razn_h_mem[15824] = 240;
razn_h_mem[15825] = 116;
razn_h_mem[15826] = 246;
razn_h_mem[15827] = 122;
razn_h_mem[15828] = 252;
razn_h_mem[15829] = 128;
razn_h_mem[15830] = 4;
razn_h_mem[15831] = 134;
razn_h_mem[15832] = 10;
razn_h_mem[15833] = 140;
razn_h_mem[15834] = 16;
razn_h_mem[15835] = 146;
razn_h_mem[15836] = 22;
razn_h_mem[15837] = 152;
razn_h_mem[15838] = 28;
razn_h_mem[15839] = 158;
razn_h_mem[15840] = 34;
razn_h_mem[15841] = 164;
razn_h_mem[15842] = 40;
razn_h_mem[15843] = 170;
razn_h_mem[15844] = 46;
razn_h_mem[15845] = 176;
razn_h_mem[15846] = 52;
razn_h_mem[15847] = 182;
razn_h_mem[15848] = 58;
razn_h_mem[15849] = 188;
razn_h_mem[15850] = 64;
razn_h_mem[15851] = 194;
razn_h_mem[15852] = 70;
razn_h_mem[15853] = 200;
razn_h_mem[15854] = 76;
razn_h_mem[15855] = 206;
razn_h_mem[15856] = 82;
razn_h_mem[15857] = 212;
razn_h_mem[15858] = 88;
razn_h_mem[15859] = 218;
razn_h_mem[15860] = 94;
razn_h_mem[15861] = 224;
razn_h_mem[15862] = 100;
razn_h_mem[15863] = 230;
razn_h_mem[15864] = 106;
razn_h_mem[15865] = 236;
razn_h_mem[15866] = 112;
razn_h_mem[15867] = 242;
razn_h_mem[15868] = 118;
razn_h_mem[15869] = 248;
razn_h_mem[15870] = 124;
razn_h_mem[15871] = 255;
razn_h_mem[15872] = 0;
razn_h_mem[15873] = 130;
razn_h_mem[15874] = 6;
razn_h_mem[15875] = 136;
razn_h_mem[15876] = 12;
razn_h_mem[15877] = 142;
razn_h_mem[15878] = 18;
razn_h_mem[15879] = 148;
razn_h_mem[15880] = 24;
razn_h_mem[15881] = 154;
razn_h_mem[15882] = 30;
razn_h_mem[15883] = 160;
razn_h_mem[15884] = 36;
razn_h_mem[15885] = 166;
razn_h_mem[15886] = 42;
razn_h_mem[15887] = 172;
razn_h_mem[15888] = 48;
razn_h_mem[15889] = 178;
razn_h_mem[15890] = 54;
razn_h_mem[15891] = 184;
razn_h_mem[15892] = 60;
razn_h_mem[15893] = 190;
razn_h_mem[15894] = 66;
razn_h_mem[15895] = 196;
razn_h_mem[15896] = 72;
razn_h_mem[15897] = 202;
razn_h_mem[15898] = 78;
razn_h_mem[15899] = 208;
razn_h_mem[15900] = 84;
razn_h_mem[15901] = 214;
razn_h_mem[15902] = 90;
razn_h_mem[15903] = 220;
razn_h_mem[15904] = 96;
razn_h_mem[15905] = 226;
razn_h_mem[15906] = 102;
razn_h_mem[15907] = 232;
razn_h_mem[15908] = 108;
razn_h_mem[15909] = 238;
razn_h_mem[15910] = 114;
razn_h_mem[15911] = 244;
razn_h_mem[15912] = 120;
razn_h_mem[15913] = 250;
razn_h_mem[15914] = 126;
razn_h_mem[15915] = 2;
razn_h_mem[15916] = 132;
razn_h_mem[15917] = 8;
razn_h_mem[15918] = 138;
razn_h_mem[15919] = 14;
razn_h_mem[15920] = 144;
razn_h_mem[15921] = 20;
razn_h_mem[15922] = 150;
razn_h_mem[15923] = 26;
razn_h_mem[15924] = 156;
razn_h_mem[15925] = 32;
razn_h_mem[15926] = 162;
razn_h_mem[15927] = 38;
razn_h_mem[15928] = 168;
razn_h_mem[15929] = 44;
razn_h_mem[15930] = 174;
razn_h_mem[15931] = 50;
razn_h_mem[15932] = 180;
razn_h_mem[15933] = 56;
razn_h_mem[15934] = 186;
razn_h_mem[15935] = 62;
razn_h_mem[15936] = 192;
razn_h_mem[15937] = 68;
razn_h_mem[15938] = 198;
razn_h_mem[15939] = 74;
razn_h_mem[15940] = 204;
razn_h_mem[15941] = 80;
razn_h_mem[15942] = 210;
razn_h_mem[15943] = 86;
razn_h_mem[15944] = 216;
razn_h_mem[15945] = 92;
razn_h_mem[15946] = 222;
razn_h_mem[15947] = 98;
razn_h_mem[15948] = 228;
razn_h_mem[15949] = 104;
razn_h_mem[15950] = 234;
razn_h_mem[15951] = 110;
razn_h_mem[15952] = 240;
razn_h_mem[15953] = 116;
razn_h_mem[15954] = 246;
razn_h_mem[15955] = 122;
razn_h_mem[15956] = 252;
razn_h_mem[15957] = 128;
razn_h_mem[15958] = 4;
razn_h_mem[15959] = 134;
razn_h_mem[15960] = 10;
razn_h_mem[15961] = 140;
razn_h_mem[15962] = 16;
razn_h_mem[15963] = 146;
razn_h_mem[15964] = 22;
razn_h_mem[15965] = 152;
razn_h_mem[15966] = 28;
razn_h_mem[15967] = 158;
razn_h_mem[15968] = 34;
razn_h_mem[15969] = 164;
razn_h_mem[15970] = 40;
razn_h_mem[15971] = 170;
razn_h_mem[15972] = 46;
razn_h_mem[15973] = 176;
razn_h_mem[15974] = 52;
razn_h_mem[15975] = 182;
razn_h_mem[15976] = 58;
razn_h_mem[15977] = 188;
razn_h_mem[15978] = 64;
razn_h_mem[15979] = 194;
razn_h_mem[15980] = 70;
razn_h_mem[15981] = 200;
razn_h_mem[15982] = 76;
razn_h_mem[15983] = 206;
razn_h_mem[15984] = 82;
razn_h_mem[15985] = 212;
razn_h_mem[15986] = 88;
razn_h_mem[15987] = 218;
razn_h_mem[15988] = 94;
razn_h_mem[15989] = 224;
razn_h_mem[15990] = 100;
razn_h_mem[15991] = 230;
razn_h_mem[15992] = 106;
razn_h_mem[15993] = 236;
razn_h_mem[15994] = 112;
razn_h_mem[15995] = 242;
razn_h_mem[15996] = 118;
razn_h_mem[15997] = 248;
razn_h_mem[15998] = 124;
razn_h_mem[15999] = 255;
razn_h_mem[16000] = 0;
razn_h_mem[16001] = 130;
razn_h_mem[16002] = 6;
razn_h_mem[16003] = 136;
razn_h_mem[16004] = 12;
razn_h_mem[16005] = 142;
razn_h_mem[16006] = 18;
razn_h_mem[16007] = 148;
razn_h_mem[16008] = 24;
razn_h_mem[16009] = 154;
razn_h_mem[16010] = 30;
razn_h_mem[16011] = 160;
razn_h_mem[16012] = 36;
razn_h_mem[16013] = 166;
razn_h_mem[16014] = 42;
razn_h_mem[16015] = 172;
razn_h_mem[16016] = 48;
razn_h_mem[16017] = 178;
razn_h_mem[16018] = 54;
razn_h_mem[16019] = 184;
razn_h_mem[16020] = 60;
razn_h_mem[16021] = 190;
razn_h_mem[16022] = 66;
razn_h_mem[16023] = 196;
razn_h_mem[16024] = 72;
razn_h_mem[16025] = 202;
razn_h_mem[16026] = 78;
razn_h_mem[16027] = 208;
razn_h_mem[16028] = 84;
razn_h_mem[16029] = 214;
razn_h_mem[16030] = 90;
razn_h_mem[16031] = 220;
razn_h_mem[16032] = 96;
razn_h_mem[16033] = 226;
razn_h_mem[16034] = 102;
razn_h_mem[16035] = 232;
razn_h_mem[16036] = 108;
razn_h_mem[16037] = 238;
razn_h_mem[16038] = 114;
razn_h_mem[16039] = 244;
razn_h_mem[16040] = 120;
razn_h_mem[16041] = 250;
razn_h_mem[16042] = 126;
razn_h_mem[16043] = 2;
razn_h_mem[16044] = 132;
razn_h_mem[16045] = 8;
razn_h_mem[16046] = 138;
razn_h_mem[16047] = 14;
razn_h_mem[16048] = 144;
razn_h_mem[16049] = 20;
razn_h_mem[16050] = 150;
razn_h_mem[16051] = 26;
razn_h_mem[16052] = 156;
razn_h_mem[16053] = 32;
razn_h_mem[16054] = 162;
razn_h_mem[16055] = 38;
razn_h_mem[16056] = 168;
razn_h_mem[16057] = 44;
razn_h_mem[16058] = 174;
razn_h_mem[16059] = 50;
razn_h_mem[16060] = 180;
razn_h_mem[16061] = 56;
razn_h_mem[16062] = 186;
razn_h_mem[16063] = 62;
razn_h_mem[16064] = 192;
razn_h_mem[16065] = 68;
razn_h_mem[16066] = 198;
razn_h_mem[16067] = 74;
razn_h_mem[16068] = 204;
razn_h_mem[16069] = 80;
razn_h_mem[16070] = 210;
razn_h_mem[16071] = 86;
razn_h_mem[16072] = 216;
razn_h_mem[16073] = 92;
razn_h_mem[16074] = 222;
razn_h_mem[16075] = 98;
razn_h_mem[16076] = 228;
razn_h_mem[16077] = 104;
razn_h_mem[16078] = 234;
razn_h_mem[16079] = 110;
razn_h_mem[16080] = 240;
razn_h_mem[16081] = 116;
razn_h_mem[16082] = 246;
razn_h_mem[16083] = 122;
razn_h_mem[16084] = 252;
razn_h_mem[16085] = 128;
razn_h_mem[16086] = 4;
razn_h_mem[16087] = 134;
razn_h_mem[16088] = 10;
razn_h_mem[16089] = 140;
razn_h_mem[16090] = 16;
razn_h_mem[16091] = 146;
razn_h_mem[16092] = 22;
razn_h_mem[16093] = 152;
razn_h_mem[16094] = 28;
razn_h_mem[16095] = 158;
razn_h_mem[16096] = 34;
razn_h_mem[16097] = 164;
razn_h_mem[16098] = 40;
razn_h_mem[16099] = 170;
razn_h_mem[16100] = 46;
razn_h_mem[16101] = 176;
razn_h_mem[16102] = 52;
razn_h_mem[16103] = 182;
razn_h_mem[16104] = 58;
razn_h_mem[16105] = 188;
razn_h_mem[16106] = 64;
razn_h_mem[16107] = 194;
razn_h_mem[16108] = 70;
razn_h_mem[16109] = 200;
razn_h_mem[16110] = 76;
razn_h_mem[16111] = 206;
razn_h_mem[16112] = 82;
razn_h_mem[16113] = 212;
razn_h_mem[16114] = 88;
razn_h_mem[16115] = 218;
razn_h_mem[16116] = 94;
razn_h_mem[16117] = 224;
razn_h_mem[16118] = 100;
razn_h_mem[16119] = 230;
razn_h_mem[16120] = 106;
razn_h_mem[16121] = 236;
razn_h_mem[16122] = 112;
razn_h_mem[16123] = 242;
razn_h_mem[16124] = 118;
razn_h_mem[16125] = 248;
razn_h_mem[16126] = 124;
razn_h_mem[16127] = 255;
razn_h_mem[16128] = 0;
razn_h_mem[16129] = 130;
razn_h_mem[16130] = 6;
razn_h_mem[16131] = 136;
razn_h_mem[16132] = 12;
razn_h_mem[16133] = 142;
razn_h_mem[16134] = 18;
razn_h_mem[16135] = 148;
razn_h_mem[16136] = 24;
razn_h_mem[16137] = 154;
razn_h_mem[16138] = 30;
razn_h_mem[16139] = 160;
razn_h_mem[16140] = 36;
razn_h_mem[16141] = 166;
razn_h_mem[16142] = 42;
razn_h_mem[16143] = 172;
razn_h_mem[16144] = 48;
razn_h_mem[16145] = 178;
razn_h_mem[16146] = 54;
razn_h_mem[16147] = 184;
razn_h_mem[16148] = 60;
razn_h_mem[16149] = 190;
razn_h_mem[16150] = 66;
razn_h_mem[16151] = 196;
razn_h_mem[16152] = 72;
razn_h_mem[16153] = 202;
razn_h_mem[16154] = 78;
razn_h_mem[16155] = 208;
razn_h_mem[16156] = 84;
razn_h_mem[16157] = 214;
razn_h_mem[16158] = 90;
razn_h_mem[16159] = 220;
razn_h_mem[16160] = 96;
razn_h_mem[16161] = 226;
razn_h_mem[16162] = 102;
razn_h_mem[16163] = 232;
razn_h_mem[16164] = 108;
razn_h_mem[16165] = 238;
razn_h_mem[16166] = 114;
razn_h_mem[16167] = 244;
razn_h_mem[16168] = 120;
razn_h_mem[16169] = 250;
razn_h_mem[16170] = 126;
razn_h_mem[16171] = 2;
razn_h_mem[16172] = 132;
razn_h_mem[16173] = 8;
razn_h_mem[16174] = 138;
razn_h_mem[16175] = 14;
razn_h_mem[16176] = 144;
razn_h_mem[16177] = 20;
razn_h_mem[16178] = 150;
razn_h_mem[16179] = 26;
razn_h_mem[16180] = 156;
razn_h_mem[16181] = 32;
razn_h_mem[16182] = 162;
razn_h_mem[16183] = 38;
razn_h_mem[16184] = 168;
razn_h_mem[16185] = 44;
razn_h_mem[16186] = 174;
razn_h_mem[16187] = 50;
razn_h_mem[16188] = 180;
razn_h_mem[16189] = 56;
razn_h_mem[16190] = 186;
razn_h_mem[16191] = 62;
razn_h_mem[16192] = 192;
razn_h_mem[16193] = 68;
razn_h_mem[16194] = 198;
razn_h_mem[16195] = 74;
razn_h_mem[16196] = 204;
razn_h_mem[16197] = 80;
razn_h_mem[16198] = 210;
razn_h_mem[16199] = 86;
razn_h_mem[16200] = 216;
razn_h_mem[16201] = 92;
razn_h_mem[16202] = 222;
razn_h_mem[16203] = 98;
razn_h_mem[16204] = 228;
razn_h_mem[16205] = 104;
razn_h_mem[16206] = 234;
razn_h_mem[16207] = 110;
razn_h_mem[16208] = 240;
razn_h_mem[16209] = 116;
razn_h_mem[16210] = 246;
razn_h_mem[16211] = 122;
razn_h_mem[16212] = 252;
razn_h_mem[16213] = 128;
razn_h_mem[16214] = 4;
razn_h_mem[16215] = 134;
razn_h_mem[16216] = 10;
razn_h_mem[16217] = 140;
razn_h_mem[16218] = 16;
razn_h_mem[16219] = 146;
razn_h_mem[16220] = 22;
razn_h_mem[16221] = 152;
razn_h_mem[16222] = 28;
razn_h_mem[16223] = 158;
razn_h_mem[16224] = 34;
razn_h_mem[16225] = 164;
razn_h_mem[16226] = 40;
razn_h_mem[16227] = 170;
razn_h_mem[16228] = 46;
razn_h_mem[16229] = 176;
razn_h_mem[16230] = 52;
razn_h_mem[16231] = 182;
razn_h_mem[16232] = 58;
razn_h_mem[16233] = 188;
razn_h_mem[16234] = 64;
razn_h_mem[16235] = 194;
razn_h_mem[16236] = 70;
razn_h_mem[16237] = 200;
razn_h_mem[16238] = 76;
razn_h_mem[16239] = 206;
razn_h_mem[16240] = 82;
razn_h_mem[16241] = 212;
razn_h_mem[16242] = 88;
razn_h_mem[16243] = 218;
razn_h_mem[16244] = 94;
razn_h_mem[16245] = 224;
razn_h_mem[16246] = 100;
razn_h_mem[16247] = 230;
razn_h_mem[16248] = 106;
razn_h_mem[16249] = 236;
razn_h_mem[16250] = 112;
razn_h_mem[16251] = 242;
razn_h_mem[16252] = 118;
razn_h_mem[16253] = 248;
razn_h_mem[16254] = 124;
razn_h_mem[16255] = 255;
razn_h_mem[16256] = 0;
razn_h_mem[16257] = 130;
razn_h_mem[16258] = 6;
razn_h_mem[16259] = 136;
razn_h_mem[16260] = 12;
razn_h_mem[16261] = 142;
razn_h_mem[16262] = 18;
razn_h_mem[16263] = 148;
razn_h_mem[16264] = 24;
razn_h_mem[16265] = 154;
razn_h_mem[16266] = 30;
razn_h_mem[16267] = 160;
razn_h_mem[16268] = 36;
razn_h_mem[16269] = 166;
razn_h_mem[16270] = 42;
razn_h_mem[16271] = 172;
razn_h_mem[16272] = 48;
razn_h_mem[16273] = 178;
razn_h_mem[16274] = 54;
razn_h_mem[16275] = 184;
razn_h_mem[16276] = 60;
razn_h_mem[16277] = 190;
razn_h_mem[16278] = 66;
razn_h_mem[16279] = 196;
razn_h_mem[16280] = 72;
razn_h_mem[16281] = 202;
razn_h_mem[16282] = 78;
razn_h_mem[16283] = 208;
razn_h_mem[16284] = 84;
razn_h_mem[16285] = 214;
razn_h_mem[16286] = 90;
razn_h_mem[16287] = 220;
razn_h_mem[16288] = 96;
razn_h_mem[16289] = 226;
razn_h_mem[16290] = 102;
razn_h_mem[16291] = 232;
razn_h_mem[16292] = 108;
razn_h_mem[16293] = 238;
razn_h_mem[16294] = 114;
razn_h_mem[16295] = 244;
razn_h_mem[16296] = 120;
razn_h_mem[16297] = 250;
razn_h_mem[16298] = 126;
razn_h_mem[16299] = 2;
razn_h_mem[16300] = 132;
razn_h_mem[16301] = 8;
razn_h_mem[16302] = 138;
razn_h_mem[16303] = 14;
razn_h_mem[16304] = 144;
razn_h_mem[16305] = 20;
razn_h_mem[16306] = 150;
razn_h_mem[16307] = 26;
razn_h_mem[16308] = 156;
razn_h_mem[16309] = 32;
razn_h_mem[16310] = 162;
razn_h_mem[16311] = 38;
razn_h_mem[16312] = 168;
razn_h_mem[16313] = 44;
razn_h_mem[16314] = 174;
razn_h_mem[16315] = 50;
razn_h_mem[16316] = 180;
razn_h_mem[16317] = 56;
razn_h_mem[16318] = 186;
razn_h_mem[16319] = 62;
razn_h_mem[16320] = 192;
razn_h_mem[16321] = 68;
razn_h_mem[16322] = 198;
razn_h_mem[16323] = 74;
razn_h_mem[16324] = 204;
razn_h_mem[16325] = 80;
razn_h_mem[16326] = 210;
razn_h_mem[16327] = 86;
razn_h_mem[16328] = 216;
razn_h_mem[16329] = 92;
razn_h_mem[16330] = 222;
razn_h_mem[16331] = 98;
razn_h_mem[16332] = 228;
razn_h_mem[16333] = 104;
razn_h_mem[16334] = 234;
razn_h_mem[16335] = 110;
razn_h_mem[16336] = 240;
razn_h_mem[16337] = 116;
razn_h_mem[16338] = 246;
razn_h_mem[16339] = 122;
razn_h_mem[16340] = 252;
razn_h_mem[16341] = 128;
razn_h_mem[16342] = 4;
razn_h_mem[16343] = 134;
razn_h_mem[16344] = 10;
razn_h_mem[16345] = 140;
razn_h_mem[16346] = 16;
razn_h_mem[16347] = 146;
razn_h_mem[16348] = 22;
razn_h_mem[16349] = 152;
razn_h_mem[16350] = 28;
razn_h_mem[16351] = 158;
razn_h_mem[16352] = 34;
razn_h_mem[16353] = 164;
razn_h_mem[16354] = 40;
razn_h_mem[16355] = 170;
razn_h_mem[16356] = 46;
razn_h_mem[16357] = 176;
razn_h_mem[16358] = 52;
razn_h_mem[16359] = 182;
razn_h_mem[16360] = 58;
razn_h_mem[16361] = 188;
razn_h_mem[16362] = 64;
razn_h_mem[16363] = 194;
razn_h_mem[16364] = 70;
razn_h_mem[16365] = 200;
razn_h_mem[16366] = 76;
razn_h_mem[16367] = 206;
razn_h_mem[16368] = 82;
razn_h_mem[16369] = 212;
razn_h_mem[16370] = 88;
razn_h_mem[16371] = 218;
razn_h_mem[16372] = 94;
razn_h_mem[16373] = 224;
razn_h_mem[16374] = 100;
razn_h_mem[16375] = 230;
razn_h_mem[16376] = 106;
razn_h_mem[16377] = 236;
razn_h_mem[16378] = 112;
razn_h_mem[16379] = 242;
razn_h_mem[16380] = 118;
razn_h_mem[16381] = 248;
razn_h_mem[16382] = 124;
razn_h_mem[16383] = 255;
end
initial
begin
razn_w_mem[0] = 0;
razn_w_mem[1] = 0;
razn_w_mem[2] = 0;
razn_w_mem[3] = 0;
razn_w_mem[4] = 0;
razn_w_mem[5] = 0;
razn_w_mem[6] = 0;
razn_w_mem[7] = 0;
razn_w_mem[8] = 0;
razn_w_mem[9] = 0;
razn_w_mem[10] = 0;
razn_w_mem[11] = 0;
razn_w_mem[12] = 0;
razn_w_mem[13] = 0;
razn_w_mem[14] = 0;
razn_w_mem[15] = 0;
razn_w_mem[16] = 0;
razn_w_mem[17] = 0;
razn_w_mem[18] = 0;
razn_w_mem[19] = 0;
razn_w_mem[20] = 0;
razn_w_mem[21] = 0;
razn_w_mem[22] = 0;
razn_w_mem[23] = 0;
razn_w_mem[24] = 0;
razn_w_mem[25] = 0;
razn_w_mem[26] = 0;
razn_w_mem[27] = 0;
razn_w_mem[28] = 0;
razn_w_mem[29] = 0;
razn_w_mem[30] = 0;
razn_w_mem[31] = 0;
razn_w_mem[32] = 0;
razn_w_mem[33] = 0;
razn_w_mem[34] = 0;
razn_w_mem[35] = 0;
razn_w_mem[36] = 0;
razn_w_mem[37] = 0;
razn_w_mem[38] = 0;
razn_w_mem[39] = 0;
razn_w_mem[40] = 0;
razn_w_mem[41] = 0;
razn_w_mem[42] = 0;
razn_w_mem[43] = 0;
razn_w_mem[44] = 0;
razn_w_mem[45] = 0;
razn_w_mem[46] = 0;
razn_w_mem[47] = 0;
razn_w_mem[48] = 0;
razn_w_mem[49] = 0;
razn_w_mem[50] = 0;
razn_w_mem[51] = 0;
razn_w_mem[52] = 0;
razn_w_mem[53] = 0;
razn_w_mem[54] = 0;
razn_w_mem[55] = 0;
razn_w_mem[56] = 0;
razn_w_mem[57] = 0;
razn_w_mem[58] = 0;
razn_w_mem[59] = 0;
razn_w_mem[60] = 0;
razn_w_mem[61] = 0;
razn_w_mem[62] = 0;
razn_w_mem[63] = 0;
razn_w_mem[64] = 0;
razn_w_mem[65] = 0;
razn_w_mem[66] = 0;
razn_w_mem[67] = 0;
razn_w_mem[68] = 0;
razn_w_mem[69] = 0;
razn_w_mem[70] = 0;
razn_w_mem[71] = 0;
razn_w_mem[72] = 0;
razn_w_mem[73] = 0;
razn_w_mem[74] = 0;
razn_w_mem[75] = 0;
razn_w_mem[76] = 0;
razn_w_mem[77] = 0;
razn_w_mem[78] = 0;
razn_w_mem[79] = 0;
razn_w_mem[80] = 0;
razn_w_mem[81] = 0;
razn_w_mem[82] = 0;
razn_w_mem[83] = 0;
razn_w_mem[84] = 0;
razn_w_mem[85] = 0;
razn_w_mem[86] = 0;
razn_w_mem[87] = 0;
razn_w_mem[88] = 0;
razn_w_mem[89] = 0;
razn_w_mem[90] = 0;
razn_w_mem[91] = 0;
razn_w_mem[92] = 0;
razn_w_mem[93] = 0;
razn_w_mem[94] = 0;
razn_w_mem[95] = 0;
razn_w_mem[96] = 0;
razn_w_mem[97] = 0;
razn_w_mem[98] = 0;
razn_w_mem[99] = 0;
razn_w_mem[100] = 0;
razn_w_mem[101] = 0;
razn_w_mem[102] = 0;
razn_w_mem[103] = 0;
razn_w_mem[104] = 0;
razn_w_mem[105] = 0;
razn_w_mem[106] = 0;
razn_w_mem[107] = 0;
razn_w_mem[108] = 0;
razn_w_mem[109] = 0;
razn_w_mem[110] = 0;
razn_w_mem[111] = 0;
razn_w_mem[112] = 0;
razn_w_mem[113] = 0;
razn_w_mem[114] = 0;
razn_w_mem[115] = 0;
razn_w_mem[116] = 0;
razn_w_mem[117] = 0;
razn_w_mem[118] = 0;
razn_w_mem[119] = 0;
razn_w_mem[120] = 0;
razn_w_mem[121] = 0;
razn_w_mem[122] = 0;
razn_w_mem[123] = 0;
razn_w_mem[124] = 0;
razn_w_mem[125] = 0;
razn_w_mem[126] = 0;
razn_w_mem[127] = 0;
razn_w_mem[128] = 224;
razn_w_mem[129] = 224;
razn_w_mem[130] = 224;
razn_w_mem[131] = 224;
razn_w_mem[132] = 224;
razn_w_mem[133] = 224;
razn_w_mem[134] = 224;
razn_w_mem[135] = 224;
razn_w_mem[136] = 224;
razn_w_mem[137] = 224;
razn_w_mem[138] = 224;
razn_w_mem[139] = 224;
razn_w_mem[140] = 224;
razn_w_mem[141] = 224;
razn_w_mem[142] = 224;
razn_w_mem[143] = 224;
razn_w_mem[144] = 224;
razn_w_mem[145] = 224;
razn_w_mem[146] = 224;
razn_w_mem[147] = 224;
razn_w_mem[148] = 224;
razn_w_mem[149] = 224;
razn_w_mem[150] = 224;
razn_w_mem[151] = 224;
razn_w_mem[152] = 224;
razn_w_mem[153] = 224;
razn_w_mem[154] = 224;
razn_w_mem[155] = 224;
razn_w_mem[156] = 224;
razn_w_mem[157] = 224;
razn_w_mem[158] = 224;
razn_w_mem[159] = 224;
razn_w_mem[160] = 224;
razn_w_mem[161] = 224;
razn_w_mem[162] = 224;
razn_w_mem[163] = 224;
razn_w_mem[164] = 224;
razn_w_mem[165] = 224;
razn_w_mem[166] = 224;
razn_w_mem[167] = 224;
razn_w_mem[168] = 224;
razn_w_mem[169] = 224;
razn_w_mem[170] = 224;
razn_w_mem[171] = 224;
razn_w_mem[172] = 224;
razn_w_mem[173] = 224;
razn_w_mem[174] = 224;
razn_w_mem[175] = 224;
razn_w_mem[176] = 224;
razn_w_mem[177] = 224;
razn_w_mem[178] = 224;
razn_w_mem[179] = 224;
razn_w_mem[180] = 224;
razn_w_mem[181] = 224;
razn_w_mem[182] = 224;
razn_w_mem[183] = 224;
razn_w_mem[184] = 224;
razn_w_mem[185] = 224;
razn_w_mem[186] = 224;
razn_w_mem[187] = 224;
razn_w_mem[188] = 224;
razn_w_mem[189] = 224;
razn_w_mem[190] = 224;
razn_w_mem[191] = 224;
razn_w_mem[192] = 224;
razn_w_mem[193] = 224;
razn_w_mem[194] = 224;
razn_w_mem[195] = 224;
razn_w_mem[196] = 224;
razn_w_mem[197] = 224;
razn_w_mem[198] = 224;
razn_w_mem[199] = 224;
razn_w_mem[200] = 224;
razn_w_mem[201] = 224;
razn_w_mem[202] = 224;
razn_w_mem[203] = 224;
razn_w_mem[204] = 224;
razn_w_mem[205] = 224;
razn_w_mem[206] = 224;
razn_w_mem[207] = 224;
razn_w_mem[208] = 224;
razn_w_mem[209] = 224;
razn_w_mem[210] = 224;
razn_w_mem[211] = 224;
razn_w_mem[212] = 224;
razn_w_mem[213] = 224;
razn_w_mem[214] = 224;
razn_w_mem[215] = 224;
razn_w_mem[216] = 224;
razn_w_mem[217] = 224;
razn_w_mem[218] = 224;
razn_w_mem[219] = 224;
razn_w_mem[220] = 224;
razn_w_mem[221] = 224;
razn_w_mem[222] = 224;
razn_w_mem[223] = 224;
razn_w_mem[224] = 224;
razn_w_mem[225] = 224;
razn_w_mem[226] = 224;
razn_w_mem[227] = 224;
razn_w_mem[228] = 224;
razn_w_mem[229] = 224;
razn_w_mem[230] = 224;
razn_w_mem[231] = 224;
razn_w_mem[232] = 224;
razn_w_mem[233] = 224;
razn_w_mem[234] = 224;
razn_w_mem[235] = 224;
razn_w_mem[236] = 224;
razn_w_mem[237] = 224;
razn_w_mem[238] = 224;
razn_w_mem[239] = 224;
razn_w_mem[240] = 224;
razn_w_mem[241] = 224;
razn_w_mem[242] = 224;
razn_w_mem[243] = 224;
razn_w_mem[244] = 224;
razn_w_mem[245] = 224;
razn_w_mem[246] = 224;
razn_w_mem[247] = 224;
razn_w_mem[248] = 224;
razn_w_mem[249] = 224;
razn_w_mem[250] = 224;
razn_w_mem[251] = 224;
razn_w_mem[252] = 224;
razn_w_mem[253] = 224;
razn_w_mem[254] = 224;
razn_w_mem[255] = 224;
razn_w_mem[256] = 194;
razn_w_mem[257] = 194;
razn_w_mem[258] = 194;
razn_w_mem[259] = 194;
razn_w_mem[260] = 194;
razn_w_mem[261] = 194;
razn_w_mem[262] = 194;
razn_w_mem[263] = 194;
razn_w_mem[264] = 194;
razn_w_mem[265] = 194;
razn_w_mem[266] = 194;
razn_w_mem[267] = 194;
razn_w_mem[268] = 194;
razn_w_mem[269] = 194;
razn_w_mem[270] = 194;
razn_w_mem[271] = 194;
razn_w_mem[272] = 194;
razn_w_mem[273] = 194;
razn_w_mem[274] = 194;
razn_w_mem[275] = 194;
razn_w_mem[276] = 194;
razn_w_mem[277] = 194;
razn_w_mem[278] = 194;
razn_w_mem[279] = 194;
razn_w_mem[280] = 194;
razn_w_mem[281] = 194;
razn_w_mem[282] = 194;
razn_w_mem[283] = 194;
razn_w_mem[284] = 194;
razn_w_mem[285] = 194;
razn_w_mem[286] = 194;
razn_w_mem[287] = 194;
razn_w_mem[288] = 194;
razn_w_mem[289] = 194;
razn_w_mem[290] = 194;
razn_w_mem[291] = 194;
razn_w_mem[292] = 194;
razn_w_mem[293] = 194;
razn_w_mem[294] = 194;
razn_w_mem[295] = 194;
razn_w_mem[296] = 194;
razn_w_mem[297] = 194;
razn_w_mem[298] = 194;
razn_w_mem[299] = 194;
razn_w_mem[300] = 194;
razn_w_mem[301] = 194;
razn_w_mem[302] = 194;
razn_w_mem[303] = 194;
razn_w_mem[304] = 194;
razn_w_mem[305] = 194;
razn_w_mem[306] = 194;
razn_w_mem[307] = 194;
razn_w_mem[308] = 194;
razn_w_mem[309] = 194;
razn_w_mem[310] = 194;
razn_w_mem[311] = 194;
razn_w_mem[312] = 194;
razn_w_mem[313] = 194;
razn_w_mem[314] = 194;
razn_w_mem[315] = 194;
razn_w_mem[316] = 194;
razn_w_mem[317] = 194;
razn_w_mem[318] = 194;
razn_w_mem[319] = 194;
razn_w_mem[320] = 194;
razn_w_mem[321] = 194;
razn_w_mem[322] = 194;
razn_w_mem[323] = 194;
razn_w_mem[324] = 194;
razn_w_mem[325] = 194;
razn_w_mem[326] = 194;
razn_w_mem[327] = 194;
razn_w_mem[328] = 194;
razn_w_mem[329] = 194;
razn_w_mem[330] = 194;
razn_w_mem[331] = 194;
razn_w_mem[332] = 194;
razn_w_mem[333] = 194;
razn_w_mem[334] = 194;
razn_w_mem[335] = 194;
razn_w_mem[336] = 194;
razn_w_mem[337] = 194;
razn_w_mem[338] = 194;
razn_w_mem[339] = 194;
razn_w_mem[340] = 194;
razn_w_mem[341] = 194;
razn_w_mem[342] = 194;
razn_w_mem[343] = 194;
razn_w_mem[344] = 194;
razn_w_mem[345] = 194;
razn_w_mem[346] = 194;
razn_w_mem[347] = 194;
razn_w_mem[348] = 194;
razn_w_mem[349] = 194;
razn_w_mem[350] = 194;
razn_w_mem[351] = 194;
razn_w_mem[352] = 194;
razn_w_mem[353] = 194;
razn_w_mem[354] = 194;
razn_w_mem[355] = 194;
razn_w_mem[356] = 194;
razn_w_mem[357] = 194;
razn_w_mem[358] = 194;
razn_w_mem[359] = 194;
razn_w_mem[360] = 194;
razn_w_mem[361] = 194;
razn_w_mem[362] = 194;
razn_w_mem[363] = 194;
razn_w_mem[364] = 194;
razn_w_mem[365] = 194;
razn_w_mem[366] = 194;
razn_w_mem[367] = 194;
razn_w_mem[368] = 194;
razn_w_mem[369] = 194;
razn_w_mem[370] = 194;
razn_w_mem[371] = 194;
razn_w_mem[372] = 194;
razn_w_mem[373] = 194;
razn_w_mem[374] = 194;
razn_w_mem[375] = 194;
razn_w_mem[376] = 194;
razn_w_mem[377] = 194;
razn_w_mem[378] = 194;
razn_w_mem[379] = 194;
razn_w_mem[380] = 194;
razn_w_mem[381] = 194;
razn_w_mem[382] = 194;
razn_w_mem[383] = 194;
razn_w_mem[384] = 164;
razn_w_mem[385] = 164;
razn_w_mem[386] = 164;
razn_w_mem[387] = 164;
razn_w_mem[388] = 164;
razn_w_mem[389] = 164;
razn_w_mem[390] = 164;
razn_w_mem[391] = 164;
razn_w_mem[392] = 164;
razn_w_mem[393] = 164;
razn_w_mem[394] = 164;
razn_w_mem[395] = 164;
razn_w_mem[396] = 164;
razn_w_mem[397] = 164;
razn_w_mem[398] = 164;
razn_w_mem[399] = 164;
razn_w_mem[400] = 164;
razn_w_mem[401] = 164;
razn_w_mem[402] = 164;
razn_w_mem[403] = 164;
razn_w_mem[404] = 164;
razn_w_mem[405] = 164;
razn_w_mem[406] = 164;
razn_w_mem[407] = 164;
razn_w_mem[408] = 164;
razn_w_mem[409] = 164;
razn_w_mem[410] = 164;
razn_w_mem[411] = 164;
razn_w_mem[412] = 164;
razn_w_mem[413] = 164;
razn_w_mem[414] = 164;
razn_w_mem[415] = 164;
razn_w_mem[416] = 164;
razn_w_mem[417] = 164;
razn_w_mem[418] = 164;
razn_w_mem[419] = 164;
razn_w_mem[420] = 164;
razn_w_mem[421] = 164;
razn_w_mem[422] = 164;
razn_w_mem[423] = 164;
razn_w_mem[424] = 164;
razn_w_mem[425] = 164;
razn_w_mem[426] = 164;
razn_w_mem[427] = 164;
razn_w_mem[428] = 164;
razn_w_mem[429] = 164;
razn_w_mem[430] = 164;
razn_w_mem[431] = 164;
razn_w_mem[432] = 164;
razn_w_mem[433] = 164;
razn_w_mem[434] = 164;
razn_w_mem[435] = 164;
razn_w_mem[436] = 164;
razn_w_mem[437] = 164;
razn_w_mem[438] = 164;
razn_w_mem[439] = 164;
razn_w_mem[440] = 164;
razn_w_mem[441] = 164;
razn_w_mem[442] = 164;
razn_w_mem[443] = 164;
razn_w_mem[444] = 164;
razn_w_mem[445] = 164;
razn_w_mem[446] = 164;
razn_w_mem[447] = 164;
razn_w_mem[448] = 164;
razn_w_mem[449] = 164;
razn_w_mem[450] = 164;
razn_w_mem[451] = 164;
razn_w_mem[452] = 164;
razn_w_mem[453] = 164;
razn_w_mem[454] = 164;
razn_w_mem[455] = 164;
razn_w_mem[456] = 164;
razn_w_mem[457] = 164;
razn_w_mem[458] = 164;
razn_w_mem[459] = 164;
razn_w_mem[460] = 164;
razn_w_mem[461] = 164;
razn_w_mem[462] = 164;
razn_w_mem[463] = 164;
razn_w_mem[464] = 164;
razn_w_mem[465] = 164;
razn_w_mem[466] = 164;
razn_w_mem[467] = 164;
razn_w_mem[468] = 164;
razn_w_mem[469] = 164;
razn_w_mem[470] = 164;
razn_w_mem[471] = 164;
razn_w_mem[472] = 164;
razn_w_mem[473] = 164;
razn_w_mem[474] = 164;
razn_w_mem[475] = 164;
razn_w_mem[476] = 164;
razn_w_mem[477] = 164;
razn_w_mem[478] = 164;
razn_w_mem[479] = 164;
razn_w_mem[480] = 164;
razn_w_mem[481] = 164;
razn_w_mem[482] = 164;
razn_w_mem[483] = 164;
razn_w_mem[484] = 164;
razn_w_mem[485] = 164;
razn_w_mem[486] = 164;
razn_w_mem[487] = 164;
razn_w_mem[488] = 164;
razn_w_mem[489] = 164;
razn_w_mem[490] = 164;
razn_w_mem[491] = 164;
razn_w_mem[492] = 164;
razn_w_mem[493] = 164;
razn_w_mem[494] = 164;
razn_w_mem[495] = 164;
razn_w_mem[496] = 164;
razn_w_mem[497] = 164;
razn_w_mem[498] = 164;
razn_w_mem[499] = 164;
razn_w_mem[500] = 164;
razn_w_mem[501] = 164;
razn_w_mem[502] = 164;
razn_w_mem[503] = 164;
razn_w_mem[504] = 164;
razn_w_mem[505] = 164;
razn_w_mem[506] = 164;
razn_w_mem[507] = 164;
razn_w_mem[508] = 164;
razn_w_mem[509] = 164;
razn_w_mem[510] = 164;
razn_w_mem[511] = 164;
razn_w_mem[512] = 134;
razn_w_mem[513] = 134;
razn_w_mem[514] = 134;
razn_w_mem[515] = 134;
razn_w_mem[516] = 134;
razn_w_mem[517] = 134;
razn_w_mem[518] = 134;
razn_w_mem[519] = 134;
razn_w_mem[520] = 134;
razn_w_mem[521] = 134;
razn_w_mem[522] = 134;
razn_w_mem[523] = 134;
razn_w_mem[524] = 134;
razn_w_mem[525] = 134;
razn_w_mem[526] = 134;
razn_w_mem[527] = 134;
razn_w_mem[528] = 134;
razn_w_mem[529] = 134;
razn_w_mem[530] = 134;
razn_w_mem[531] = 134;
razn_w_mem[532] = 134;
razn_w_mem[533] = 134;
razn_w_mem[534] = 134;
razn_w_mem[535] = 134;
razn_w_mem[536] = 134;
razn_w_mem[537] = 134;
razn_w_mem[538] = 134;
razn_w_mem[539] = 134;
razn_w_mem[540] = 134;
razn_w_mem[541] = 134;
razn_w_mem[542] = 134;
razn_w_mem[543] = 134;
razn_w_mem[544] = 134;
razn_w_mem[545] = 134;
razn_w_mem[546] = 134;
razn_w_mem[547] = 134;
razn_w_mem[548] = 134;
razn_w_mem[549] = 134;
razn_w_mem[550] = 134;
razn_w_mem[551] = 134;
razn_w_mem[552] = 134;
razn_w_mem[553] = 134;
razn_w_mem[554] = 134;
razn_w_mem[555] = 134;
razn_w_mem[556] = 134;
razn_w_mem[557] = 134;
razn_w_mem[558] = 134;
razn_w_mem[559] = 134;
razn_w_mem[560] = 134;
razn_w_mem[561] = 134;
razn_w_mem[562] = 134;
razn_w_mem[563] = 134;
razn_w_mem[564] = 134;
razn_w_mem[565] = 134;
razn_w_mem[566] = 134;
razn_w_mem[567] = 134;
razn_w_mem[568] = 134;
razn_w_mem[569] = 134;
razn_w_mem[570] = 134;
razn_w_mem[571] = 134;
razn_w_mem[572] = 134;
razn_w_mem[573] = 134;
razn_w_mem[574] = 134;
razn_w_mem[575] = 134;
razn_w_mem[576] = 134;
razn_w_mem[577] = 134;
razn_w_mem[578] = 134;
razn_w_mem[579] = 134;
razn_w_mem[580] = 134;
razn_w_mem[581] = 134;
razn_w_mem[582] = 134;
razn_w_mem[583] = 134;
razn_w_mem[584] = 134;
razn_w_mem[585] = 134;
razn_w_mem[586] = 134;
razn_w_mem[587] = 134;
razn_w_mem[588] = 134;
razn_w_mem[589] = 134;
razn_w_mem[590] = 134;
razn_w_mem[591] = 134;
razn_w_mem[592] = 134;
razn_w_mem[593] = 134;
razn_w_mem[594] = 134;
razn_w_mem[595] = 134;
razn_w_mem[596] = 134;
razn_w_mem[597] = 134;
razn_w_mem[598] = 134;
razn_w_mem[599] = 134;
razn_w_mem[600] = 134;
razn_w_mem[601] = 134;
razn_w_mem[602] = 134;
razn_w_mem[603] = 134;
razn_w_mem[604] = 134;
razn_w_mem[605] = 134;
razn_w_mem[606] = 134;
razn_w_mem[607] = 134;
razn_w_mem[608] = 134;
razn_w_mem[609] = 134;
razn_w_mem[610] = 134;
razn_w_mem[611] = 134;
razn_w_mem[612] = 134;
razn_w_mem[613] = 134;
razn_w_mem[614] = 134;
razn_w_mem[615] = 134;
razn_w_mem[616] = 134;
razn_w_mem[617] = 134;
razn_w_mem[618] = 134;
razn_w_mem[619] = 134;
razn_w_mem[620] = 134;
razn_w_mem[621] = 134;
razn_w_mem[622] = 134;
razn_w_mem[623] = 134;
razn_w_mem[624] = 134;
razn_w_mem[625] = 134;
razn_w_mem[626] = 134;
razn_w_mem[627] = 134;
razn_w_mem[628] = 134;
razn_w_mem[629] = 134;
razn_w_mem[630] = 134;
razn_w_mem[631] = 134;
razn_w_mem[632] = 134;
razn_w_mem[633] = 134;
razn_w_mem[634] = 134;
razn_w_mem[635] = 134;
razn_w_mem[636] = 134;
razn_w_mem[637] = 134;
razn_w_mem[638] = 134;
razn_w_mem[639] = 134;
razn_w_mem[640] = 104;
razn_w_mem[641] = 104;
razn_w_mem[642] = 104;
razn_w_mem[643] = 104;
razn_w_mem[644] = 104;
razn_w_mem[645] = 104;
razn_w_mem[646] = 104;
razn_w_mem[647] = 104;
razn_w_mem[648] = 104;
razn_w_mem[649] = 104;
razn_w_mem[650] = 104;
razn_w_mem[651] = 104;
razn_w_mem[652] = 104;
razn_w_mem[653] = 104;
razn_w_mem[654] = 104;
razn_w_mem[655] = 104;
razn_w_mem[656] = 104;
razn_w_mem[657] = 104;
razn_w_mem[658] = 104;
razn_w_mem[659] = 104;
razn_w_mem[660] = 104;
razn_w_mem[661] = 104;
razn_w_mem[662] = 104;
razn_w_mem[663] = 104;
razn_w_mem[664] = 104;
razn_w_mem[665] = 104;
razn_w_mem[666] = 104;
razn_w_mem[667] = 104;
razn_w_mem[668] = 104;
razn_w_mem[669] = 104;
razn_w_mem[670] = 104;
razn_w_mem[671] = 104;
razn_w_mem[672] = 104;
razn_w_mem[673] = 104;
razn_w_mem[674] = 104;
razn_w_mem[675] = 104;
razn_w_mem[676] = 104;
razn_w_mem[677] = 104;
razn_w_mem[678] = 104;
razn_w_mem[679] = 104;
razn_w_mem[680] = 104;
razn_w_mem[681] = 104;
razn_w_mem[682] = 104;
razn_w_mem[683] = 104;
razn_w_mem[684] = 104;
razn_w_mem[685] = 104;
razn_w_mem[686] = 104;
razn_w_mem[687] = 104;
razn_w_mem[688] = 104;
razn_w_mem[689] = 104;
razn_w_mem[690] = 104;
razn_w_mem[691] = 104;
razn_w_mem[692] = 104;
razn_w_mem[693] = 104;
razn_w_mem[694] = 104;
razn_w_mem[695] = 104;
razn_w_mem[696] = 104;
razn_w_mem[697] = 104;
razn_w_mem[698] = 104;
razn_w_mem[699] = 104;
razn_w_mem[700] = 104;
razn_w_mem[701] = 104;
razn_w_mem[702] = 104;
razn_w_mem[703] = 104;
razn_w_mem[704] = 104;
razn_w_mem[705] = 104;
razn_w_mem[706] = 104;
razn_w_mem[707] = 104;
razn_w_mem[708] = 104;
razn_w_mem[709] = 104;
razn_w_mem[710] = 104;
razn_w_mem[711] = 104;
razn_w_mem[712] = 104;
razn_w_mem[713] = 104;
razn_w_mem[714] = 104;
razn_w_mem[715] = 104;
razn_w_mem[716] = 104;
razn_w_mem[717] = 104;
razn_w_mem[718] = 104;
razn_w_mem[719] = 104;
razn_w_mem[720] = 104;
razn_w_mem[721] = 104;
razn_w_mem[722] = 104;
razn_w_mem[723] = 104;
razn_w_mem[724] = 104;
razn_w_mem[725] = 104;
razn_w_mem[726] = 104;
razn_w_mem[727] = 104;
razn_w_mem[728] = 104;
razn_w_mem[729] = 104;
razn_w_mem[730] = 104;
razn_w_mem[731] = 104;
razn_w_mem[732] = 104;
razn_w_mem[733] = 104;
razn_w_mem[734] = 104;
razn_w_mem[735] = 104;
razn_w_mem[736] = 104;
razn_w_mem[737] = 104;
razn_w_mem[738] = 104;
razn_w_mem[739] = 104;
razn_w_mem[740] = 104;
razn_w_mem[741] = 104;
razn_w_mem[742] = 104;
razn_w_mem[743] = 104;
razn_w_mem[744] = 104;
razn_w_mem[745] = 104;
razn_w_mem[746] = 104;
razn_w_mem[747] = 104;
razn_w_mem[748] = 104;
razn_w_mem[749] = 104;
razn_w_mem[750] = 104;
razn_w_mem[751] = 104;
razn_w_mem[752] = 104;
razn_w_mem[753] = 104;
razn_w_mem[754] = 104;
razn_w_mem[755] = 104;
razn_w_mem[756] = 104;
razn_w_mem[757] = 104;
razn_w_mem[758] = 104;
razn_w_mem[759] = 104;
razn_w_mem[760] = 104;
razn_w_mem[761] = 104;
razn_w_mem[762] = 104;
razn_w_mem[763] = 104;
razn_w_mem[764] = 104;
razn_w_mem[765] = 104;
razn_w_mem[766] = 104;
razn_w_mem[767] = 104;
razn_w_mem[768] = 74;
razn_w_mem[769] = 74;
razn_w_mem[770] = 74;
razn_w_mem[771] = 74;
razn_w_mem[772] = 74;
razn_w_mem[773] = 74;
razn_w_mem[774] = 74;
razn_w_mem[775] = 74;
razn_w_mem[776] = 74;
razn_w_mem[777] = 74;
razn_w_mem[778] = 74;
razn_w_mem[779] = 74;
razn_w_mem[780] = 74;
razn_w_mem[781] = 74;
razn_w_mem[782] = 74;
razn_w_mem[783] = 74;
razn_w_mem[784] = 74;
razn_w_mem[785] = 74;
razn_w_mem[786] = 74;
razn_w_mem[787] = 74;
razn_w_mem[788] = 74;
razn_w_mem[789] = 74;
razn_w_mem[790] = 74;
razn_w_mem[791] = 74;
razn_w_mem[792] = 74;
razn_w_mem[793] = 74;
razn_w_mem[794] = 74;
razn_w_mem[795] = 74;
razn_w_mem[796] = 74;
razn_w_mem[797] = 74;
razn_w_mem[798] = 74;
razn_w_mem[799] = 74;
razn_w_mem[800] = 74;
razn_w_mem[801] = 74;
razn_w_mem[802] = 74;
razn_w_mem[803] = 74;
razn_w_mem[804] = 74;
razn_w_mem[805] = 74;
razn_w_mem[806] = 74;
razn_w_mem[807] = 74;
razn_w_mem[808] = 74;
razn_w_mem[809] = 74;
razn_w_mem[810] = 74;
razn_w_mem[811] = 74;
razn_w_mem[812] = 74;
razn_w_mem[813] = 74;
razn_w_mem[814] = 74;
razn_w_mem[815] = 74;
razn_w_mem[816] = 74;
razn_w_mem[817] = 74;
razn_w_mem[818] = 74;
razn_w_mem[819] = 74;
razn_w_mem[820] = 74;
razn_w_mem[821] = 74;
razn_w_mem[822] = 74;
razn_w_mem[823] = 74;
razn_w_mem[824] = 74;
razn_w_mem[825] = 74;
razn_w_mem[826] = 74;
razn_w_mem[827] = 74;
razn_w_mem[828] = 74;
razn_w_mem[829] = 74;
razn_w_mem[830] = 74;
razn_w_mem[831] = 74;
razn_w_mem[832] = 74;
razn_w_mem[833] = 74;
razn_w_mem[834] = 74;
razn_w_mem[835] = 74;
razn_w_mem[836] = 74;
razn_w_mem[837] = 74;
razn_w_mem[838] = 74;
razn_w_mem[839] = 74;
razn_w_mem[840] = 74;
razn_w_mem[841] = 74;
razn_w_mem[842] = 74;
razn_w_mem[843] = 74;
razn_w_mem[844] = 74;
razn_w_mem[845] = 74;
razn_w_mem[846] = 74;
razn_w_mem[847] = 74;
razn_w_mem[848] = 74;
razn_w_mem[849] = 74;
razn_w_mem[850] = 74;
razn_w_mem[851] = 74;
razn_w_mem[852] = 74;
razn_w_mem[853] = 74;
razn_w_mem[854] = 74;
razn_w_mem[855] = 74;
razn_w_mem[856] = 74;
razn_w_mem[857] = 74;
razn_w_mem[858] = 74;
razn_w_mem[859] = 74;
razn_w_mem[860] = 74;
razn_w_mem[861] = 74;
razn_w_mem[862] = 74;
razn_w_mem[863] = 74;
razn_w_mem[864] = 74;
razn_w_mem[865] = 74;
razn_w_mem[866] = 74;
razn_w_mem[867] = 74;
razn_w_mem[868] = 74;
razn_w_mem[869] = 74;
razn_w_mem[870] = 74;
razn_w_mem[871] = 74;
razn_w_mem[872] = 74;
razn_w_mem[873] = 74;
razn_w_mem[874] = 74;
razn_w_mem[875] = 74;
razn_w_mem[876] = 74;
razn_w_mem[877] = 74;
razn_w_mem[878] = 74;
razn_w_mem[879] = 74;
razn_w_mem[880] = 74;
razn_w_mem[881] = 74;
razn_w_mem[882] = 74;
razn_w_mem[883] = 74;
razn_w_mem[884] = 74;
razn_w_mem[885] = 74;
razn_w_mem[886] = 74;
razn_w_mem[887] = 74;
razn_w_mem[888] = 74;
razn_w_mem[889] = 74;
razn_w_mem[890] = 74;
razn_w_mem[891] = 74;
razn_w_mem[892] = 74;
razn_w_mem[893] = 74;
razn_w_mem[894] = 74;
razn_w_mem[895] = 74;
razn_w_mem[896] = 44;
razn_w_mem[897] = 44;
razn_w_mem[898] = 44;
razn_w_mem[899] = 44;
razn_w_mem[900] = 44;
razn_w_mem[901] = 44;
razn_w_mem[902] = 44;
razn_w_mem[903] = 44;
razn_w_mem[904] = 44;
razn_w_mem[905] = 44;
razn_w_mem[906] = 44;
razn_w_mem[907] = 44;
razn_w_mem[908] = 44;
razn_w_mem[909] = 44;
razn_w_mem[910] = 44;
razn_w_mem[911] = 44;
razn_w_mem[912] = 44;
razn_w_mem[913] = 44;
razn_w_mem[914] = 44;
razn_w_mem[915] = 44;
razn_w_mem[916] = 44;
razn_w_mem[917] = 44;
razn_w_mem[918] = 44;
razn_w_mem[919] = 44;
razn_w_mem[920] = 44;
razn_w_mem[921] = 44;
razn_w_mem[922] = 44;
razn_w_mem[923] = 44;
razn_w_mem[924] = 44;
razn_w_mem[925] = 44;
razn_w_mem[926] = 44;
razn_w_mem[927] = 44;
razn_w_mem[928] = 44;
razn_w_mem[929] = 44;
razn_w_mem[930] = 44;
razn_w_mem[931] = 44;
razn_w_mem[932] = 44;
razn_w_mem[933] = 44;
razn_w_mem[934] = 44;
razn_w_mem[935] = 44;
razn_w_mem[936] = 44;
razn_w_mem[937] = 44;
razn_w_mem[938] = 44;
razn_w_mem[939] = 44;
razn_w_mem[940] = 44;
razn_w_mem[941] = 44;
razn_w_mem[942] = 44;
razn_w_mem[943] = 44;
razn_w_mem[944] = 44;
razn_w_mem[945] = 44;
razn_w_mem[946] = 44;
razn_w_mem[947] = 44;
razn_w_mem[948] = 44;
razn_w_mem[949] = 44;
razn_w_mem[950] = 44;
razn_w_mem[951] = 44;
razn_w_mem[952] = 44;
razn_w_mem[953] = 44;
razn_w_mem[954] = 44;
razn_w_mem[955] = 44;
razn_w_mem[956] = 44;
razn_w_mem[957] = 44;
razn_w_mem[958] = 44;
razn_w_mem[959] = 44;
razn_w_mem[960] = 44;
razn_w_mem[961] = 44;
razn_w_mem[962] = 44;
razn_w_mem[963] = 44;
razn_w_mem[964] = 44;
razn_w_mem[965] = 44;
razn_w_mem[966] = 44;
razn_w_mem[967] = 44;
razn_w_mem[968] = 44;
razn_w_mem[969] = 44;
razn_w_mem[970] = 44;
razn_w_mem[971] = 44;
razn_w_mem[972] = 44;
razn_w_mem[973] = 44;
razn_w_mem[974] = 44;
razn_w_mem[975] = 44;
razn_w_mem[976] = 44;
razn_w_mem[977] = 44;
razn_w_mem[978] = 44;
razn_w_mem[979] = 44;
razn_w_mem[980] = 44;
razn_w_mem[981] = 44;
razn_w_mem[982] = 44;
razn_w_mem[983] = 44;
razn_w_mem[984] = 44;
razn_w_mem[985] = 44;
razn_w_mem[986] = 44;
razn_w_mem[987] = 44;
razn_w_mem[988] = 44;
razn_w_mem[989] = 44;
razn_w_mem[990] = 44;
razn_w_mem[991] = 44;
razn_w_mem[992] = 44;
razn_w_mem[993] = 44;
razn_w_mem[994] = 44;
razn_w_mem[995] = 44;
razn_w_mem[996] = 44;
razn_w_mem[997] = 44;
razn_w_mem[998] = 44;
razn_w_mem[999] = 44;
razn_w_mem[1000] = 44;
razn_w_mem[1001] = 44;
razn_w_mem[1002] = 44;
razn_w_mem[1003] = 44;
razn_w_mem[1004] = 44;
razn_w_mem[1005] = 44;
razn_w_mem[1006] = 44;
razn_w_mem[1007] = 44;
razn_w_mem[1008] = 44;
razn_w_mem[1009] = 44;
razn_w_mem[1010] = 44;
razn_w_mem[1011] = 44;
razn_w_mem[1012] = 44;
razn_w_mem[1013] = 44;
razn_w_mem[1014] = 44;
razn_w_mem[1015] = 44;
razn_w_mem[1016] = 44;
razn_w_mem[1017] = 44;
razn_w_mem[1018] = 44;
razn_w_mem[1019] = 44;
razn_w_mem[1020] = 44;
razn_w_mem[1021] = 44;
razn_w_mem[1022] = 44;
razn_w_mem[1023] = 44;
razn_w_mem[1024] = 14;
razn_w_mem[1025] = 14;
razn_w_mem[1026] = 14;
razn_w_mem[1027] = 14;
razn_w_mem[1028] = 14;
razn_w_mem[1029] = 14;
razn_w_mem[1030] = 14;
razn_w_mem[1031] = 14;
razn_w_mem[1032] = 14;
razn_w_mem[1033] = 14;
razn_w_mem[1034] = 14;
razn_w_mem[1035] = 14;
razn_w_mem[1036] = 14;
razn_w_mem[1037] = 14;
razn_w_mem[1038] = 14;
razn_w_mem[1039] = 14;
razn_w_mem[1040] = 14;
razn_w_mem[1041] = 14;
razn_w_mem[1042] = 14;
razn_w_mem[1043] = 14;
razn_w_mem[1044] = 14;
razn_w_mem[1045] = 14;
razn_w_mem[1046] = 14;
razn_w_mem[1047] = 14;
razn_w_mem[1048] = 14;
razn_w_mem[1049] = 14;
razn_w_mem[1050] = 14;
razn_w_mem[1051] = 14;
razn_w_mem[1052] = 14;
razn_w_mem[1053] = 14;
razn_w_mem[1054] = 14;
razn_w_mem[1055] = 14;
razn_w_mem[1056] = 14;
razn_w_mem[1057] = 14;
razn_w_mem[1058] = 14;
razn_w_mem[1059] = 14;
razn_w_mem[1060] = 14;
razn_w_mem[1061] = 14;
razn_w_mem[1062] = 14;
razn_w_mem[1063] = 14;
razn_w_mem[1064] = 14;
razn_w_mem[1065] = 14;
razn_w_mem[1066] = 14;
razn_w_mem[1067] = 14;
razn_w_mem[1068] = 14;
razn_w_mem[1069] = 14;
razn_w_mem[1070] = 14;
razn_w_mem[1071] = 14;
razn_w_mem[1072] = 14;
razn_w_mem[1073] = 14;
razn_w_mem[1074] = 14;
razn_w_mem[1075] = 14;
razn_w_mem[1076] = 14;
razn_w_mem[1077] = 14;
razn_w_mem[1078] = 14;
razn_w_mem[1079] = 14;
razn_w_mem[1080] = 14;
razn_w_mem[1081] = 14;
razn_w_mem[1082] = 14;
razn_w_mem[1083] = 14;
razn_w_mem[1084] = 14;
razn_w_mem[1085] = 14;
razn_w_mem[1086] = 14;
razn_w_mem[1087] = 14;
razn_w_mem[1088] = 14;
razn_w_mem[1089] = 14;
razn_w_mem[1090] = 14;
razn_w_mem[1091] = 14;
razn_w_mem[1092] = 14;
razn_w_mem[1093] = 14;
razn_w_mem[1094] = 14;
razn_w_mem[1095] = 14;
razn_w_mem[1096] = 14;
razn_w_mem[1097] = 14;
razn_w_mem[1098] = 14;
razn_w_mem[1099] = 14;
razn_w_mem[1100] = 14;
razn_w_mem[1101] = 14;
razn_w_mem[1102] = 14;
razn_w_mem[1103] = 14;
razn_w_mem[1104] = 14;
razn_w_mem[1105] = 14;
razn_w_mem[1106] = 14;
razn_w_mem[1107] = 14;
razn_w_mem[1108] = 14;
razn_w_mem[1109] = 14;
razn_w_mem[1110] = 14;
razn_w_mem[1111] = 14;
razn_w_mem[1112] = 14;
razn_w_mem[1113] = 14;
razn_w_mem[1114] = 14;
razn_w_mem[1115] = 14;
razn_w_mem[1116] = 14;
razn_w_mem[1117] = 14;
razn_w_mem[1118] = 14;
razn_w_mem[1119] = 14;
razn_w_mem[1120] = 14;
razn_w_mem[1121] = 14;
razn_w_mem[1122] = 14;
razn_w_mem[1123] = 14;
razn_w_mem[1124] = 14;
razn_w_mem[1125] = 14;
razn_w_mem[1126] = 14;
razn_w_mem[1127] = 14;
razn_w_mem[1128] = 14;
razn_w_mem[1129] = 14;
razn_w_mem[1130] = 14;
razn_w_mem[1131] = 14;
razn_w_mem[1132] = 14;
razn_w_mem[1133] = 14;
razn_w_mem[1134] = 14;
razn_w_mem[1135] = 14;
razn_w_mem[1136] = 14;
razn_w_mem[1137] = 14;
razn_w_mem[1138] = 14;
razn_w_mem[1139] = 14;
razn_w_mem[1140] = 14;
razn_w_mem[1141] = 14;
razn_w_mem[1142] = 14;
razn_w_mem[1143] = 14;
razn_w_mem[1144] = 14;
razn_w_mem[1145] = 14;
razn_w_mem[1146] = 14;
razn_w_mem[1147] = 14;
razn_w_mem[1148] = 14;
razn_w_mem[1149] = 14;
razn_w_mem[1150] = 14;
razn_w_mem[1151] = 14;
razn_w_mem[1152] = 238;
razn_w_mem[1153] = 238;
razn_w_mem[1154] = 238;
razn_w_mem[1155] = 238;
razn_w_mem[1156] = 238;
razn_w_mem[1157] = 238;
razn_w_mem[1158] = 238;
razn_w_mem[1159] = 238;
razn_w_mem[1160] = 238;
razn_w_mem[1161] = 238;
razn_w_mem[1162] = 238;
razn_w_mem[1163] = 238;
razn_w_mem[1164] = 238;
razn_w_mem[1165] = 238;
razn_w_mem[1166] = 238;
razn_w_mem[1167] = 238;
razn_w_mem[1168] = 238;
razn_w_mem[1169] = 238;
razn_w_mem[1170] = 238;
razn_w_mem[1171] = 238;
razn_w_mem[1172] = 238;
razn_w_mem[1173] = 238;
razn_w_mem[1174] = 238;
razn_w_mem[1175] = 238;
razn_w_mem[1176] = 238;
razn_w_mem[1177] = 238;
razn_w_mem[1178] = 238;
razn_w_mem[1179] = 238;
razn_w_mem[1180] = 238;
razn_w_mem[1181] = 238;
razn_w_mem[1182] = 238;
razn_w_mem[1183] = 238;
razn_w_mem[1184] = 238;
razn_w_mem[1185] = 238;
razn_w_mem[1186] = 238;
razn_w_mem[1187] = 238;
razn_w_mem[1188] = 238;
razn_w_mem[1189] = 238;
razn_w_mem[1190] = 238;
razn_w_mem[1191] = 238;
razn_w_mem[1192] = 238;
razn_w_mem[1193] = 238;
razn_w_mem[1194] = 238;
razn_w_mem[1195] = 238;
razn_w_mem[1196] = 238;
razn_w_mem[1197] = 238;
razn_w_mem[1198] = 238;
razn_w_mem[1199] = 238;
razn_w_mem[1200] = 238;
razn_w_mem[1201] = 238;
razn_w_mem[1202] = 238;
razn_w_mem[1203] = 238;
razn_w_mem[1204] = 238;
razn_w_mem[1205] = 238;
razn_w_mem[1206] = 238;
razn_w_mem[1207] = 238;
razn_w_mem[1208] = 238;
razn_w_mem[1209] = 238;
razn_w_mem[1210] = 238;
razn_w_mem[1211] = 238;
razn_w_mem[1212] = 238;
razn_w_mem[1213] = 238;
razn_w_mem[1214] = 238;
razn_w_mem[1215] = 238;
razn_w_mem[1216] = 238;
razn_w_mem[1217] = 238;
razn_w_mem[1218] = 238;
razn_w_mem[1219] = 238;
razn_w_mem[1220] = 238;
razn_w_mem[1221] = 238;
razn_w_mem[1222] = 238;
razn_w_mem[1223] = 238;
razn_w_mem[1224] = 238;
razn_w_mem[1225] = 238;
razn_w_mem[1226] = 238;
razn_w_mem[1227] = 238;
razn_w_mem[1228] = 238;
razn_w_mem[1229] = 238;
razn_w_mem[1230] = 238;
razn_w_mem[1231] = 238;
razn_w_mem[1232] = 238;
razn_w_mem[1233] = 238;
razn_w_mem[1234] = 238;
razn_w_mem[1235] = 238;
razn_w_mem[1236] = 238;
razn_w_mem[1237] = 238;
razn_w_mem[1238] = 238;
razn_w_mem[1239] = 238;
razn_w_mem[1240] = 238;
razn_w_mem[1241] = 238;
razn_w_mem[1242] = 238;
razn_w_mem[1243] = 238;
razn_w_mem[1244] = 238;
razn_w_mem[1245] = 238;
razn_w_mem[1246] = 238;
razn_w_mem[1247] = 238;
razn_w_mem[1248] = 238;
razn_w_mem[1249] = 238;
razn_w_mem[1250] = 238;
razn_w_mem[1251] = 238;
razn_w_mem[1252] = 238;
razn_w_mem[1253] = 238;
razn_w_mem[1254] = 238;
razn_w_mem[1255] = 238;
razn_w_mem[1256] = 238;
razn_w_mem[1257] = 238;
razn_w_mem[1258] = 238;
razn_w_mem[1259] = 238;
razn_w_mem[1260] = 238;
razn_w_mem[1261] = 238;
razn_w_mem[1262] = 238;
razn_w_mem[1263] = 238;
razn_w_mem[1264] = 238;
razn_w_mem[1265] = 238;
razn_w_mem[1266] = 238;
razn_w_mem[1267] = 238;
razn_w_mem[1268] = 238;
razn_w_mem[1269] = 238;
razn_w_mem[1270] = 238;
razn_w_mem[1271] = 238;
razn_w_mem[1272] = 238;
razn_w_mem[1273] = 238;
razn_w_mem[1274] = 238;
razn_w_mem[1275] = 238;
razn_w_mem[1276] = 238;
razn_w_mem[1277] = 238;
razn_w_mem[1278] = 238;
razn_w_mem[1279] = 238;
razn_w_mem[1280] = 208;
razn_w_mem[1281] = 208;
razn_w_mem[1282] = 208;
razn_w_mem[1283] = 208;
razn_w_mem[1284] = 208;
razn_w_mem[1285] = 208;
razn_w_mem[1286] = 208;
razn_w_mem[1287] = 208;
razn_w_mem[1288] = 208;
razn_w_mem[1289] = 208;
razn_w_mem[1290] = 208;
razn_w_mem[1291] = 208;
razn_w_mem[1292] = 208;
razn_w_mem[1293] = 208;
razn_w_mem[1294] = 208;
razn_w_mem[1295] = 208;
razn_w_mem[1296] = 208;
razn_w_mem[1297] = 208;
razn_w_mem[1298] = 208;
razn_w_mem[1299] = 208;
razn_w_mem[1300] = 208;
razn_w_mem[1301] = 208;
razn_w_mem[1302] = 208;
razn_w_mem[1303] = 208;
razn_w_mem[1304] = 208;
razn_w_mem[1305] = 208;
razn_w_mem[1306] = 208;
razn_w_mem[1307] = 208;
razn_w_mem[1308] = 208;
razn_w_mem[1309] = 208;
razn_w_mem[1310] = 208;
razn_w_mem[1311] = 208;
razn_w_mem[1312] = 208;
razn_w_mem[1313] = 208;
razn_w_mem[1314] = 208;
razn_w_mem[1315] = 208;
razn_w_mem[1316] = 208;
razn_w_mem[1317] = 208;
razn_w_mem[1318] = 208;
razn_w_mem[1319] = 208;
razn_w_mem[1320] = 208;
razn_w_mem[1321] = 208;
razn_w_mem[1322] = 208;
razn_w_mem[1323] = 208;
razn_w_mem[1324] = 208;
razn_w_mem[1325] = 208;
razn_w_mem[1326] = 208;
razn_w_mem[1327] = 208;
razn_w_mem[1328] = 208;
razn_w_mem[1329] = 208;
razn_w_mem[1330] = 208;
razn_w_mem[1331] = 208;
razn_w_mem[1332] = 208;
razn_w_mem[1333] = 208;
razn_w_mem[1334] = 208;
razn_w_mem[1335] = 208;
razn_w_mem[1336] = 208;
razn_w_mem[1337] = 208;
razn_w_mem[1338] = 208;
razn_w_mem[1339] = 208;
razn_w_mem[1340] = 208;
razn_w_mem[1341] = 208;
razn_w_mem[1342] = 208;
razn_w_mem[1343] = 208;
razn_w_mem[1344] = 208;
razn_w_mem[1345] = 208;
razn_w_mem[1346] = 208;
razn_w_mem[1347] = 208;
razn_w_mem[1348] = 208;
razn_w_mem[1349] = 208;
razn_w_mem[1350] = 208;
razn_w_mem[1351] = 208;
razn_w_mem[1352] = 208;
razn_w_mem[1353] = 208;
razn_w_mem[1354] = 208;
razn_w_mem[1355] = 208;
razn_w_mem[1356] = 208;
razn_w_mem[1357] = 208;
razn_w_mem[1358] = 208;
razn_w_mem[1359] = 208;
razn_w_mem[1360] = 208;
razn_w_mem[1361] = 208;
razn_w_mem[1362] = 208;
razn_w_mem[1363] = 208;
razn_w_mem[1364] = 208;
razn_w_mem[1365] = 208;
razn_w_mem[1366] = 208;
razn_w_mem[1367] = 208;
razn_w_mem[1368] = 208;
razn_w_mem[1369] = 208;
razn_w_mem[1370] = 208;
razn_w_mem[1371] = 208;
razn_w_mem[1372] = 208;
razn_w_mem[1373] = 208;
razn_w_mem[1374] = 208;
razn_w_mem[1375] = 208;
razn_w_mem[1376] = 208;
razn_w_mem[1377] = 208;
razn_w_mem[1378] = 208;
razn_w_mem[1379] = 208;
razn_w_mem[1380] = 208;
razn_w_mem[1381] = 208;
razn_w_mem[1382] = 208;
razn_w_mem[1383] = 208;
razn_w_mem[1384] = 208;
razn_w_mem[1385] = 208;
razn_w_mem[1386] = 208;
razn_w_mem[1387] = 208;
razn_w_mem[1388] = 208;
razn_w_mem[1389] = 208;
razn_w_mem[1390] = 208;
razn_w_mem[1391] = 208;
razn_w_mem[1392] = 208;
razn_w_mem[1393] = 208;
razn_w_mem[1394] = 208;
razn_w_mem[1395] = 208;
razn_w_mem[1396] = 208;
razn_w_mem[1397] = 208;
razn_w_mem[1398] = 208;
razn_w_mem[1399] = 208;
razn_w_mem[1400] = 208;
razn_w_mem[1401] = 208;
razn_w_mem[1402] = 208;
razn_w_mem[1403] = 208;
razn_w_mem[1404] = 208;
razn_w_mem[1405] = 208;
razn_w_mem[1406] = 208;
razn_w_mem[1407] = 208;
razn_w_mem[1408] = 178;
razn_w_mem[1409] = 178;
razn_w_mem[1410] = 178;
razn_w_mem[1411] = 178;
razn_w_mem[1412] = 178;
razn_w_mem[1413] = 178;
razn_w_mem[1414] = 178;
razn_w_mem[1415] = 178;
razn_w_mem[1416] = 178;
razn_w_mem[1417] = 178;
razn_w_mem[1418] = 178;
razn_w_mem[1419] = 178;
razn_w_mem[1420] = 178;
razn_w_mem[1421] = 178;
razn_w_mem[1422] = 178;
razn_w_mem[1423] = 178;
razn_w_mem[1424] = 178;
razn_w_mem[1425] = 178;
razn_w_mem[1426] = 178;
razn_w_mem[1427] = 178;
razn_w_mem[1428] = 178;
razn_w_mem[1429] = 178;
razn_w_mem[1430] = 178;
razn_w_mem[1431] = 178;
razn_w_mem[1432] = 178;
razn_w_mem[1433] = 178;
razn_w_mem[1434] = 178;
razn_w_mem[1435] = 178;
razn_w_mem[1436] = 178;
razn_w_mem[1437] = 178;
razn_w_mem[1438] = 178;
razn_w_mem[1439] = 178;
razn_w_mem[1440] = 178;
razn_w_mem[1441] = 178;
razn_w_mem[1442] = 178;
razn_w_mem[1443] = 178;
razn_w_mem[1444] = 178;
razn_w_mem[1445] = 178;
razn_w_mem[1446] = 178;
razn_w_mem[1447] = 178;
razn_w_mem[1448] = 178;
razn_w_mem[1449] = 178;
razn_w_mem[1450] = 178;
razn_w_mem[1451] = 178;
razn_w_mem[1452] = 178;
razn_w_mem[1453] = 178;
razn_w_mem[1454] = 178;
razn_w_mem[1455] = 178;
razn_w_mem[1456] = 178;
razn_w_mem[1457] = 178;
razn_w_mem[1458] = 178;
razn_w_mem[1459] = 178;
razn_w_mem[1460] = 178;
razn_w_mem[1461] = 178;
razn_w_mem[1462] = 178;
razn_w_mem[1463] = 178;
razn_w_mem[1464] = 178;
razn_w_mem[1465] = 178;
razn_w_mem[1466] = 178;
razn_w_mem[1467] = 178;
razn_w_mem[1468] = 178;
razn_w_mem[1469] = 178;
razn_w_mem[1470] = 178;
razn_w_mem[1471] = 178;
razn_w_mem[1472] = 178;
razn_w_mem[1473] = 178;
razn_w_mem[1474] = 178;
razn_w_mem[1475] = 178;
razn_w_mem[1476] = 178;
razn_w_mem[1477] = 178;
razn_w_mem[1478] = 178;
razn_w_mem[1479] = 178;
razn_w_mem[1480] = 178;
razn_w_mem[1481] = 178;
razn_w_mem[1482] = 178;
razn_w_mem[1483] = 178;
razn_w_mem[1484] = 178;
razn_w_mem[1485] = 178;
razn_w_mem[1486] = 178;
razn_w_mem[1487] = 178;
razn_w_mem[1488] = 178;
razn_w_mem[1489] = 178;
razn_w_mem[1490] = 178;
razn_w_mem[1491] = 178;
razn_w_mem[1492] = 178;
razn_w_mem[1493] = 178;
razn_w_mem[1494] = 178;
razn_w_mem[1495] = 178;
razn_w_mem[1496] = 178;
razn_w_mem[1497] = 178;
razn_w_mem[1498] = 178;
razn_w_mem[1499] = 178;
razn_w_mem[1500] = 178;
razn_w_mem[1501] = 178;
razn_w_mem[1502] = 178;
razn_w_mem[1503] = 178;
razn_w_mem[1504] = 178;
razn_w_mem[1505] = 178;
razn_w_mem[1506] = 178;
razn_w_mem[1507] = 178;
razn_w_mem[1508] = 178;
razn_w_mem[1509] = 178;
razn_w_mem[1510] = 178;
razn_w_mem[1511] = 178;
razn_w_mem[1512] = 178;
razn_w_mem[1513] = 178;
razn_w_mem[1514] = 178;
razn_w_mem[1515] = 178;
razn_w_mem[1516] = 178;
razn_w_mem[1517] = 178;
razn_w_mem[1518] = 178;
razn_w_mem[1519] = 178;
razn_w_mem[1520] = 178;
razn_w_mem[1521] = 178;
razn_w_mem[1522] = 178;
razn_w_mem[1523] = 178;
razn_w_mem[1524] = 178;
razn_w_mem[1525] = 178;
razn_w_mem[1526] = 178;
razn_w_mem[1527] = 178;
razn_w_mem[1528] = 178;
razn_w_mem[1529] = 178;
razn_w_mem[1530] = 178;
razn_w_mem[1531] = 178;
razn_w_mem[1532] = 178;
razn_w_mem[1533] = 178;
razn_w_mem[1534] = 178;
razn_w_mem[1535] = 178;
razn_w_mem[1536] = 148;
razn_w_mem[1537] = 148;
razn_w_mem[1538] = 148;
razn_w_mem[1539] = 148;
razn_w_mem[1540] = 148;
razn_w_mem[1541] = 148;
razn_w_mem[1542] = 148;
razn_w_mem[1543] = 148;
razn_w_mem[1544] = 148;
razn_w_mem[1545] = 148;
razn_w_mem[1546] = 148;
razn_w_mem[1547] = 148;
razn_w_mem[1548] = 148;
razn_w_mem[1549] = 148;
razn_w_mem[1550] = 148;
razn_w_mem[1551] = 148;
razn_w_mem[1552] = 148;
razn_w_mem[1553] = 148;
razn_w_mem[1554] = 148;
razn_w_mem[1555] = 148;
razn_w_mem[1556] = 148;
razn_w_mem[1557] = 148;
razn_w_mem[1558] = 148;
razn_w_mem[1559] = 148;
razn_w_mem[1560] = 148;
razn_w_mem[1561] = 148;
razn_w_mem[1562] = 148;
razn_w_mem[1563] = 148;
razn_w_mem[1564] = 148;
razn_w_mem[1565] = 148;
razn_w_mem[1566] = 148;
razn_w_mem[1567] = 148;
razn_w_mem[1568] = 148;
razn_w_mem[1569] = 148;
razn_w_mem[1570] = 148;
razn_w_mem[1571] = 148;
razn_w_mem[1572] = 148;
razn_w_mem[1573] = 148;
razn_w_mem[1574] = 148;
razn_w_mem[1575] = 148;
razn_w_mem[1576] = 148;
razn_w_mem[1577] = 148;
razn_w_mem[1578] = 148;
razn_w_mem[1579] = 148;
razn_w_mem[1580] = 148;
razn_w_mem[1581] = 148;
razn_w_mem[1582] = 148;
razn_w_mem[1583] = 148;
razn_w_mem[1584] = 148;
razn_w_mem[1585] = 148;
razn_w_mem[1586] = 148;
razn_w_mem[1587] = 148;
razn_w_mem[1588] = 148;
razn_w_mem[1589] = 148;
razn_w_mem[1590] = 148;
razn_w_mem[1591] = 148;
razn_w_mem[1592] = 148;
razn_w_mem[1593] = 148;
razn_w_mem[1594] = 148;
razn_w_mem[1595] = 148;
razn_w_mem[1596] = 148;
razn_w_mem[1597] = 148;
razn_w_mem[1598] = 148;
razn_w_mem[1599] = 148;
razn_w_mem[1600] = 148;
razn_w_mem[1601] = 148;
razn_w_mem[1602] = 148;
razn_w_mem[1603] = 148;
razn_w_mem[1604] = 148;
razn_w_mem[1605] = 148;
razn_w_mem[1606] = 148;
razn_w_mem[1607] = 148;
razn_w_mem[1608] = 148;
razn_w_mem[1609] = 148;
razn_w_mem[1610] = 148;
razn_w_mem[1611] = 148;
razn_w_mem[1612] = 148;
razn_w_mem[1613] = 148;
razn_w_mem[1614] = 148;
razn_w_mem[1615] = 148;
razn_w_mem[1616] = 148;
razn_w_mem[1617] = 148;
razn_w_mem[1618] = 148;
razn_w_mem[1619] = 148;
razn_w_mem[1620] = 148;
razn_w_mem[1621] = 148;
razn_w_mem[1622] = 148;
razn_w_mem[1623] = 148;
razn_w_mem[1624] = 148;
razn_w_mem[1625] = 148;
razn_w_mem[1626] = 148;
razn_w_mem[1627] = 148;
razn_w_mem[1628] = 148;
razn_w_mem[1629] = 148;
razn_w_mem[1630] = 148;
razn_w_mem[1631] = 148;
razn_w_mem[1632] = 148;
razn_w_mem[1633] = 148;
razn_w_mem[1634] = 148;
razn_w_mem[1635] = 148;
razn_w_mem[1636] = 148;
razn_w_mem[1637] = 148;
razn_w_mem[1638] = 148;
razn_w_mem[1639] = 148;
razn_w_mem[1640] = 148;
razn_w_mem[1641] = 148;
razn_w_mem[1642] = 148;
razn_w_mem[1643] = 148;
razn_w_mem[1644] = 148;
razn_w_mem[1645] = 148;
razn_w_mem[1646] = 148;
razn_w_mem[1647] = 148;
razn_w_mem[1648] = 148;
razn_w_mem[1649] = 148;
razn_w_mem[1650] = 148;
razn_w_mem[1651] = 148;
razn_w_mem[1652] = 148;
razn_w_mem[1653] = 148;
razn_w_mem[1654] = 148;
razn_w_mem[1655] = 148;
razn_w_mem[1656] = 148;
razn_w_mem[1657] = 148;
razn_w_mem[1658] = 148;
razn_w_mem[1659] = 148;
razn_w_mem[1660] = 148;
razn_w_mem[1661] = 148;
razn_w_mem[1662] = 148;
razn_w_mem[1663] = 148;
razn_w_mem[1664] = 118;
razn_w_mem[1665] = 118;
razn_w_mem[1666] = 118;
razn_w_mem[1667] = 118;
razn_w_mem[1668] = 118;
razn_w_mem[1669] = 118;
razn_w_mem[1670] = 118;
razn_w_mem[1671] = 118;
razn_w_mem[1672] = 118;
razn_w_mem[1673] = 118;
razn_w_mem[1674] = 118;
razn_w_mem[1675] = 118;
razn_w_mem[1676] = 118;
razn_w_mem[1677] = 118;
razn_w_mem[1678] = 118;
razn_w_mem[1679] = 118;
razn_w_mem[1680] = 118;
razn_w_mem[1681] = 118;
razn_w_mem[1682] = 118;
razn_w_mem[1683] = 118;
razn_w_mem[1684] = 118;
razn_w_mem[1685] = 118;
razn_w_mem[1686] = 118;
razn_w_mem[1687] = 118;
razn_w_mem[1688] = 118;
razn_w_mem[1689] = 118;
razn_w_mem[1690] = 118;
razn_w_mem[1691] = 118;
razn_w_mem[1692] = 118;
razn_w_mem[1693] = 118;
razn_w_mem[1694] = 118;
razn_w_mem[1695] = 118;
razn_w_mem[1696] = 118;
razn_w_mem[1697] = 118;
razn_w_mem[1698] = 118;
razn_w_mem[1699] = 118;
razn_w_mem[1700] = 118;
razn_w_mem[1701] = 118;
razn_w_mem[1702] = 118;
razn_w_mem[1703] = 118;
razn_w_mem[1704] = 118;
razn_w_mem[1705] = 118;
razn_w_mem[1706] = 118;
razn_w_mem[1707] = 118;
razn_w_mem[1708] = 118;
razn_w_mem[1709] = 118;
razn_w_mem[1710] = 118;
razn_w_mem[1711] = 118;
razn_w_mem[1712] = 118;
razn_w_mem[1713] = 118;
razn_w_mem[1714] = 118;
razn_w_mem[1715] = 118;
razn_w_mem[1716] = 118;
razn_w_mem[1717] = 118;
razn_w_mem[1718] = 118;
razn_w_mem[1719] = 118;
razn_w_mem[1720] = 118;
razn_w_mem[1721] = 118;
razn_w_mem[1722] = 118;
razn_w_mem[1723] = 118;
razn_w_mem[1724] = 118;
razn_w_mem[1725] = 118;
razn_w_mem[1726] = 118;
razn_w_mem[1727] = 118;
razn_w_mem[1728] = 118;
razn_w_mem[1729] = 118;
razn_w_mem[1730] = 118;
razn_w_mem[1731] = 118;
razn_w_mem[1732] = 118;
razn_w_mem[1733] = 118;
razn_w_mem[1734] = 118;
razn_w_mem[1735] = 118;
razn_w_mem[1736] = 118;
razn_w_mem[1737] = 118;
razn_w_mem[1738] = 118;
razn_w_mem[1739] = 118;
razn_w_mem[1740] = 118;
razn_w_mem[1741] = 118;
razn_w_mem[1742] = 118;
razn_w_mem[1743] = 118;
razn_w_mem[1744] = 118;
razn_w_mem[1745] = 118;
razn_w_mem[1746] = 118;
razn_w_mem[1747] = 118;
razn_w_mem[1748] = 118;
razn_w_mem[1749] = 118;
razn_w_mem[1750] = 118;
razn_w_mem[1751] = 118;
razn_w_mem[1752] = 118;
razn_w_mem[1753] = 118;
razn_w_mem[1754] = 118;
razn_w_mem[1755] = 118;
razn_w_mem[1756] = 118;
razn_w_mem[1757] = 118;
razn_w_mem[1758] = 118;
razn_w_mem[1759] = 118;
razn_w_mem[1760] = 118;
razn_w_mem[1761] = 118;
razn_w_mem[1762] = 118;
razn_w_mem[1763] = 118;
razn_w_mem[1764] = 118;
razn_w_mem[1765] = 118;
razn_w_mem[1766] = 118;
razn_w_mem[1767] = 118;
razn_w_mem[1768] = 118;
razn_w_mem[1769] = 118;
razn_w_mem[1770] = 118;
razn_w_mem[1771] = 118;
razn_w_mem[1772] = 118;
razn_w_mem[1773] = 118;
razn_w_mem[1774] = 118;
razn_w_mem[1775] = 118;
razn_w_mem[1776] = 118;
razn_w_mem[1777] = 118;
razn_w_mem[1778] = 118;
razn_w_mem[1779] = 118;
razn_w_mem[1780] = 118;
razn_w_mem[1781] = 118;
razn_w_mem[1782] = 118;
razn_w_mem[1783] = 118;
razn_w_mem[1784] = 118;
razn_w_mem[1785] = 118;
razn_w_mem[1786] = 118;
razn_w_mem[1787] = 118;
razn_w_mem[1788] = 118;
razn_w_mem[1789] = 118;
razn_w_mem[1790] = 118;
razn_w_mem[1791] = 118;
razn_w_mem[1792] = 88;
razn_w_mem[1793] = 88;
razn_w_mem[1794] = 88;
razn_w_mem[1795] = 88;
razn_w_mem[1796] = 88;
razn_w_mem[1797] = 88;
razn_w_mem[1798] = 88;
razn_w_mem[1799] = 88;
razn_w_mem[1800] = 88;
razn_w_mem[1801] = 88;
razn_w_mem[1802] = 88;
razn_w_mem[1803] = 88;
razn_w_mem[1804] = 88;
razn_w_mem[1805] = 88;
razn_w_mem[1806] = 88;
razn_w_mem[1807] = 88;
razn_w_mem[1808] = 88;
razn_w_mem[1809] = 88;
razn_w_mem[1810] = 88;
razn_w_mem[1811] = 88;
razn_w_mem[1812] = 88;
razn_w_mem[1813] = 88;
razn_w_mem[1814] = 88;
razn_w_mem[1815] = 88;
razn_w_mem[1816] = 88;
razn_w_mem[1817] = 88;
razn_w_mem[1818] = 88;
razn_w_mem[1819] = 88;
razn_w_mem[1820] = 88;
razn_w_mem[1821] = 88;
razn_w_mem[1822] = 88;
razn_w_mem[1823] = 88;
razn_w_mem[1824] = 88;
razn_w_mem[1825] = 88;
razn_w_mem[1826] = 88;
razn_w_mem[1827] = 88;
razn_w_mem[1828] = 88;
razn_w_mem[1829] = 88;
razn_w_mem[1830] = 88;
razn_w_mem[1831] = 88;
razn_w_mem[1832] = 88;
razn_w_mem[1833] = 88;
razn_w_mem[1834] = 88;
razn_w_mem[1835] = 88;
razn_w_mem[1836] = 88;
razn_w_mem[1837] = 88;
razn_w_mem[1838] = 88;
razn_w_mem[1839] = 88;
razn_w_mem[1840] = 88;
razn_w_mem[1841] = 88;
razn_w_mem[1842] = 88;
razn_w_mem[1843] = 88;
razn_w_mem[1844] = 88;
razn_w_mem[1845] = 88;
razn_w_mem[1846] = 88;
razn_w_mem[1847] = 88;
razn_w_mem[1848] = 88;
razn_w_mem[1849] = 88;
razn_w_mem[1850] = 88;
razn_w_mem[1851] = 88;
razn_w_mem[1852] = 88;
razn_w_mem[1853] = 88;
razn_w_mem[1854] = 88;
razn_w_mem[1855] = 88;
razn_w_mem[1856] = 88;
razn_w_mem[1857] = 88;
razn_w_mem[1858] = 88;
razn_w_mem[1859] = 88;
razn_w_mem[1860] = 88;
razn_w_mem[1861] = 88;
razn_w_mem[1862] = 88;
razn_w_mem[1863] = 88;
razn_w_mem[1864] = 88;
razn_w_mem[1865] = 88;
razn_w_mem[1866] = 88;
razn_w_mem[1867] = 88;
razn_w_mem[1868] = 88;
razn_w_mem[1869] = 88;
razn_w_mem[1870] = 88;
razn_w_mem[1871] = 88;
razn_w_mem[1872] = 88;
razn_w_mem[1873] = 88;
razn_w_mem[1874] = 88;
razn_w_mem[1875] = 88;
razn_w_mem[1876] = 88;
razn_w_mem[1877] = 88;
razn_w_mem[1878] = 88;
razn_w_mem[1879] = 88;
razn_w_mem[1880] = 88;
razn_w_mem[1881] = 88;
razn_w_mem[1882] = 88;
razn_w_mem[1883] = 88;
razn_w_mem[1884] = 88;
razn_w_mem[1885] = 88;
razn_w_mem[1886] = 88;
razn_w_mem[1887] = 88;
razn_w_mem[1888] = 88;
razn_w_mem[1889] = 88;
razn_w_mem[1890] = 88;
razn_w_mem[1891] = 88;
razn_w_mem[1892] = 88;
razn_w_mem[1893] = 88;
razn_w_mem[1894] = 88;
razn_w_mem[1895] = 88;
razn_w_mem[1896] = 88;
razn_w_mem[1897] = 88;
razn_w_mem[1898] = 88;
razn_w_mem[1899] = 88;
razn_w_mem[1900] = 88;
razn_w_mem[1901] = 88;
razn_w_mem[1902] = 88;
razn_w_mem[1903] = 88;
razn_w_mem[1904] = 88;
razn_w_mem[1905] = 88;
razn_w_mem[1906] = 88;
razn_w_mem[1907] = 88;
razn_w_mem[1908] = 88;
razn_w_mem[1909] = 88;
razn_w_mem[1910] = 88;
razn_w_mem[1911] = 88;
razn_w_mem[1912] = 88;
razn_w_mem[1913] = 88;
razn_w_mem[1914] = 88;
razn_w_mem[1915] = 88;
razn_w_mem[1916] = 88;
razn_w_mem[1917] = 88;
razn_w_mem[1918] = 88;
razn_w_mem[1919] = 88;
razn_w_mem[1920] = 58;
razn_w_mem[1921] = 58;
razn_w_mem[1922] = 58;
razn_w_mem[1923] = 58;
razn_w_mem[1924] = 58;
razn_w_mem[1925] = 58;
razn_w_mem[1926] = 58;
razn_w_mem[1927] = 58;
razn_w_mem[1928] = 58;
razn_w_mem[1929] = 58;
razn_w_mem[1930] = 58;
razn_w_mem[1931] = 58;
razn_w_mem[1932] = 58;
razn_w_mem[1933] = 58;
razn_w_mem[1934] = 58;
razn_w_mem[1935] = 58;
razn_w_mem[1936] = 58;
razn_w_mem[1937] = 58;
razn_w_mem[1938] = 58;
razn_w_mem[1939] = 58;
razn_w_mem[1940] = 58;
razn_w_mem[1941] = 58;
razn_w_mem[1942] = 58;
razn_w_mem[1943] = 58;
razn_w_mem[1944] = 58;
razn_w_mem[1945] = 58;
razn_w_mem[1946] = 58;
razn_w_mem[1947] = 58;
razn_w_mem[1948] = 58;
razn_w_mem[1949] = 58;
razn_w_mem[1950] = 58;
razn_w_mem[1951] = 58;
razn_w_mem[1952] = 58;
razn_w_mem[1953] = 58;
razn_w_mem[1954] = 58;
razn_w_mem[1955] = 58;
razn_w_mem[1956] = 58;
razn_w_mem[1957] = 58;
razn_w_mem[1958] = 58;
razn_w_mem[1959] = 58;
razn_w_mem[1960] = 58;
razn_w_mem[1961] = 58;
razn_w_mem[1962] = 58;
razn_w_mem[1963] = 58;
razn_w_mem[1964] = 58;
razn_w_mem[1965] = 58;
razn_w_mem[1966] = 58;
razn_w_mem[1967] = 58;
razn_w_mem[1968] = 58;
razn_w_mem[1969] = 58;
razn_w_mem[1970] = 58;
razn_w_mem[1971] = 58;
razn_w_mem[1972] = 58;
razn_w_mem[1973] = 58;
razn_w_mem[1974] = 58;
razn_w_mem[1975] = 58;
razn_w_mem[1976] = 58;
razn_w_mem[1977] = 58;
razn_w_mem[1978] = 58;
razn_w_mem[1979] = 58;
razn_w_mem[1980] = 58;
razn_w_mem[1981] = 58;
razn_w_mem[1982] = 58;
razn_w_mem[1983] = 58;
razn_w_mem[1984] = 58;
razn_w_mem[1985] = 58;
razn_w_mem[1986] = 58;
razn_w_mem[1987] = 58;
razn_w_mem[1988] = 58;
razn_w_mem[1989] = 58;
razn_w_mem[1990] = 58;
razn_w_mem[1991] = 58;
razn_w_mem[1992] = 58;
razn_w_mem[1993] = 58;
razn_w_mem[1994] = 58;
razn_w_mem[1995] = 58;
razn_w_mem[1996] = 58;
razn_w_mem[1997] = 58;
razn_w_mem[1998] = 58;
razn_w_mem[1999] = 58;
razn_w_mem[2000] = 58;
razn_w_mem[2001] = 58;
razn_w_mem[2002] = 58;
razn_w_mem[2003] = 58;
razn_w_mem[2004] = 58;
razn_w_mem[2005] = 58;
razn_w_mem[2006] = 58;
razn_w_mem[2007] = 58;
razn_w_mem[2008] = 58;
razn_w_mem[2009] = 58;
razn_w_mem[2010] = 58;
razn_w_mem[2011] = 58;
razn_w_mem[2012] = 58;
razn_w_mem[2013] = 58;
razn_w_mem[2014] = 58;
razn_w_mem[2015] = 58;
razn_w_mem[2016] = 58;
razn_w_mem[2017] = 58;
razn_w_mem[2018] = 58;
razn_w_mem[2019] = 58;
razn_w_mem[2020] = 58;
razn_w_mem[2021] = 58;
razn_w_mem[2022] = 58;
razn_w_mem[2023] = 58;
razn_w_mem[2024] = 58;
razn_w_mem[2025] = 58;
razn_w_mem[2026] = 58;
razn_w_mem[2027] = 58;
razn_w_mem[2028] = 58;
razn_w_mem[2029] = 58;
razn_w_mem[2030] = 58;
razn_w_mem[2031] = 58;
razn_w_mem[2032] = 58;
razn_w_mem[2033] = 58;
razn_w_mem[2034] = 58;
razn_w_mem[2035] = 58;
razn_w_mem[2036] = 58;
razn_w_mem[2037] = 58;
razn_w_mem[2038] = 58;
razn_w_mem[2039] = 58;
razn_w_mem[2040] = 58;
razn_w_mem[2041] = 58;
razn_w_mem[2042] = 58;
razn_w_mem[2043] = 58;
razn_w_mem[2044] = 58;
razn_w_mem[2045] = 58;
razn_w_mem[2046] = 58;
razn_w_mem[2047] = 58;
razn_w_mem[2048] = 28;
razn_w_mem[2049] = 28;
razn_w_mem[2050] = 28;
razn_w_mem[2051] = 28;
razn_w_mem[2052] = 28;
razn_w_mem[2053] = 28;
razn_w_mem[2054] = 28;
razn_w_mem[2055] = 28;
razn_w_mem[2056] = 28;
razn_w_mem[2057] = 28;
razn_w_mem[2058] = 28;
razn_w_mem[2059] = 28;
razn_w_mem[2060] = 28;
razn_w_mem[2061] = 28;
razn_w_mem[2062] = 28;
razn_w_mem[2063] = 28;
razn_w_mem[2064] = 28;
razn_w_mem[2065] = 28;
razn_w_mem[2066] = 28;
razn_w_mem[2067] = 28;
razn_w_mem[2068] = 28;
razn_w_mem[2069] = 28;
razn_w_mem[2070] = 28;
razn_w_mem[2071] = 28;
razn_w_mem[2072] = 28;
razn_w_mem[2073] = 28;
razn_w_mem[2074] = 28;
razn_w_mem[2075] = 28;
razn_w_mem[2076] = 28;
razn_w_mem[2077] = 28;
razn_w_mem[2078] = 28;
razn_w_mem[2079] = 28;
razn_w_mem[2080] = 28;
razn_w_mem[2081] = 28;
razn_w_mem[2082] = 28;
razn_w_mem[2083] = 28;
razn_w_mem[2084] = 28;
razn_w_mem[2085] = 28;
razn_w_mem[2086] = 28;
razn_w_mem[2087] = 28;
razn_w_mem[2088] = 28;
razn_w_mem[2089] = 28;
razn_w_mem[2090] = 28;
razn_w_mem[2091] = 28;
razn_w_mem[2092] = 28;
razn_w_mem[2093] = 28;
razn_w_mem[2094] = 28;
razn_w_mem[2095] = 28;
razn_w_mem[2096] = 28;
razn_w_mem[2097] = 28;
razn_w_mem[2098] = 28;
razn_w_mem[2099] = 28;
razn_w_mem[2100] = 28;
razn_w_mem[2101] = 28;
razn_w_mem[2102] = 28;
razn_w_mem[2103] = 28;
razn_w_mem[2104] = 28;
razn_w_mem[2105] = 28;
razn_w_mem[2106] = 28;
razn_w_mem[2107] = 28;
razn_w_mem[2108] = 28;
razn_w_mem[2109] = 28;
razn_w_mem[2110] = 28;
razn_w_mem[2111] = 28;
razn_w_mem[2112] = 28;
razn_w_mem[2113] = 28;
razn_w_mem[2114] = 28;
razn_w_mem[2115] = 28;
razn_w_mem[2116] = 28;
razn_w_mem[2117] = 28;
razn_w_mem[2118] = 28;
razn_w_mem[2119] = 28;
razn_w_mem[2120] = 28;
razn_w_mem[2121] = 28;
razn_w_mem[2122] = 28;
razn_w_mem[2123] = 28;
razn_w_mem[2124] = 28;
razn_w_mem[2125] = 28;
razn_w_mem[2126] = 28;
razn_w_mem[2127] = 28;
razn_w_mem[2128] = 28;
razn_w_mem[2129] = 28;
razn_w_mem[2130] = 28;
razn_w_mem[2131] = 28;
razn_w_mem[2132] = 28;
razn_w_mem[2133] = 28;
razn_w_mem[2134] = 28;
razn_w_mem[2135] = 28;
razn_w_mem[2136] = 28;
razn_w_mem[2137] = 28;
razn_w_mem[2138] = 28;
razn_w_mem[2139] = 28;
razn_w_mem[2140] = 28;
razn_w_mem[2141] = 28;
razn_w_mem[2142] = 28;
razn_w_mem[2143] = 28;
razn_w_mem[2144] = 28;
razn_w_mem[2145] = 28;
razn_w_mem[2146] = 28;
razn_w_mem[2147] = 28;
razn_w_mem[2148] = 28;
razn_w_mem[2149] = 28;
razn_w_mem[2150] = 28;
razn_w_mem[2151] = 28;
razn_w_mem[2152] = 28;
razn_w_mem[2153] = 28;
razn_w_mem[2154] = 28;
razn_w_mem[2155] = 28;
razn_w_mem[2156] = 28;
razn_w_mem[2157] = 28;
razn_w_mem[2158] = 28;
razn_w_mem[2159] = 28;
razn_w_mem[2160] = 28;
razn_w_mem[2161] = 28;
razn_w_mem[2162] = 28;
razn_w_mem[2163] = 28;
razn_w_mem[2164] = 28;
razn_w_mem[2165] = 28;
razn_w_mem[2166] = 28;
razn_w_mem[2167] = 28;
razn_w_mem[2168] = 28;
razn_w_mem[2169] = 28;
razn_w_mem[2170] = 28;
razn_w_mem[2171] = 28;
razn_w_mem[2172] = 28;
razn_w_mem[2173] = 28;
razn_w_mem[2174] = 28;
razn_w_mem[2175] = 28;
razn_w_mem[2176] = 252;
razn_w_mem[2177] = 252;
razn_w_mem[2178] = 252;
razn_w_mem[2179] = 252;
razn_w_mem[2180] = 252;
razn_w_mem[2181] = 252;
razn_w_mem[2182] = 252;
razn_w_mem[2183] = 252;
razn_w_mem[2184] = 252;
razn_w_mem[2185] = 252;
razn_w_mem[2186] = 252;
razn_w_mem[2187] = 252;
razn_w_mem[2188] = 252;
razn_w_mem[2189] = 252;
razn_w_mem[2190] = 252;
razn_w_mem[2191] = 252;
razn_w_mem[2192] = 252;
razn_w_mem[2193] = 252;
razn_w_mem[2194] = 252;
razn_w_mem[2195] = 252;
razn_w_mem[2196] = 252;
razn_w_mem[2197] = 252;
razn_w_mem[2198] = 252;
razn_w_mem[2199] = 252;
razn_w_mem[2200] = 252;
razn_w_mem[2201] = 252;
razn_w_mem[2202] = 252;
razn_w_mem[2203] = 252;
razn_w_mem[2204] = 252;
razn_w_mem[2205] = 252;
razn_w_mem[2206] = 252;
razn_w_mem[2207] = 252;
razn_w_mem[2208] = 252;
razn_w_mem[2209] = 252;
razn_w_mem[2210] = 252;
razn_w_mem[2211] = 252;
razn_w_mem[2212] = 252;
razn_w_mem[2213] = 252;
razn_w_mem[2214] = 252;
razn_w_mem[2215] = 252;
razn_w_mem[2216] = 252;
razn_w_mem[2217] = 252;
razn_w_mem[2218] = 252;
razn_w_mem[2219] = 252;
razn_w_mem[2220] = 252;
razn_w_mem[2221] = 252;
razn_w_mem[2222] = 252;
razn_w_mem[2223] = 252;
razn_w_mem[2224] = 252;
razn_w_mem[2225] = 252;
razn_w_mem[2226] = 252;
razn_w_mem[2227] = 252;
razn_w_mem[2228] = 252;
razn_w_mem[2229] = 252;
razn_w_mem[2230] = 252;
razn_w_mem[2231] = 252;
razn_w_mem[2232] = 252;
razn_w_mem[2233] = 252;
razn_w_mem[2234] = 252;
razn_w_mem[2235] = 252;
razn_w_mem[2236] = 252;
razn_w_mem[2237] = 252;
razn_w_mem[2238] = 252;
razn_w_mem[2239] = 252;
razn_w_mem[2240] = 252;
razn_w_mem[2241] = 252;
razn_w_mem[2242] = 252;
razn_w_mem[2243] = 252;
razn_w_mem[2244] = 252;
razn_w_mem[2245] = 252;
razn_w_mem[2246] = 252;
razn_w_mem[2247] = 252;
razn_w_mem[2248] = 252;
razn_w_mem[2249] = 252;
razn_w_mem[2250] = 252;
razn_w_mem[2251] = 252;
razn_w_mem[2252] = 252;
razn_w_mem[2253] = 252;
razn_w_mem[2254] = 252;
razn_w_mem[2255] = 252;
razn_w_mem[2256] = 252;
razn_w_mem[2257] = 252;
razn_w_mem[2258] = 252;
razn_w_mem[2259] = 252;
razn_w_mem[2260] = 252;
razn_w_mem[2261] = 252;
razn_w_mem[2262] = 252;
razn_w_mem[2263] = 252;
razn_w_mem[2264] = 252;
razn_w_mem[2265] = 252;
razn_w_mem[2266] = 252;
razn_w_mem[2267] = 252;
razn_w_mem[2268] = 252;
razn_w_mem[2269] = 252;
razn_w_mem[2270] = 252;
razn_w_mem[2271] = 252;
razn_w_mem[2272] = 252;
razn_w_mem[2273] = 252;
razn_w_mem[2274] = 252;
razn_w_mem[2275] = 252;
razn_w_mem[2276] = 252;
razn_w_mem[2277] = 252;
razn_w_mem[2278] = 252;
razn_w_mem[2279] = 252;
razn_w_mem[2280] = 252;
razn_w_mem[2281] = 252;
razn_w_mem[2282] = 252;
razn_w_mem[2283] = 252;
razn_w_mem[2284] = 252;
razn_w_mem[2285] = 252;
razn_w_mem[2286] = 252;
razn_w_mem[2287] = 252;
razn_w_mem[2288] = 252;
razn_w_mem[2289] = 252;
razn_w_mem[2290] = 252;
razn_w_mem[2291] = 252;
razn_w_mem[2292] = 252;
razn_w_mem[2293] = 252;
razn_w_mem[2294] = 252;
razn_w_mem[2295] = 252;
razn_w_mem[2296] = 252;
razn_w_mem[2297] = 252;
razn_w_mem[2298] = 252;
razn_w_mem[2299] = 252;
razn_w_mem[2300] = 252;
razn_w_mem[2301] = 252;
razn_w_mem[2302] = 252;
razn_w_mem[2303] = 252;
razn_w_mem[2304] = 222;
razn_w_mem[2305] = 222;
razn_w_mem[2306] = 222;
razn_w_mem[2307] = 222;
razn_w_mem[2308] = 222;
razn_w_mem[2309] = 222;
razn_w_mem[2310] = 222;
razn_w_mem[2311] = 222;
razn_w_mem[2312] = 222;
razn_w_mem[2313] = 222;
razn_w_mem[2314] = 222;
razn_w_mem[2315] = 222;
razn_w_mem[2316] = 222;
razn_w_mem[2317] = 222;
razn_w_mem[2318] = 222;
razn_w_mem[2319] = 222;
razn_w_mem[2320] = 222;
razn_w_mem[2321] = 222;
razn_w_mem[2322] = 222;
razn_w_mem[2323] = 222;
razn_w_mem[2324] = 222;
razn_w_mem[2325] = 222;
razn_w_mem[2326] = 222;
razn_w_mem[2327] = 222;
razn_w_mem[2328] = 222;
razn_w_mem[2329] = 222;
razn_w_mem[2330] = 222;
razn_w_mem[2331] = 222;
razn_w_mem[2332] = 222;
razn_w_mem[2333] = 222;
razn_w_mem[2334] = 222;
razn_w_mem[2335] = 222;
razn_w_mem[2336] = 222;
razn_w_mem[2337] = 222;
razn_w_mem[2338] = 222;
razn_w_mem[2339] = 222;
razn_w_mem[2340] = 222;
razn_w_mem[2341] = 222;
razn_w_mem[2342] = 222;
razn_w_mem[2343] = 222;
razn_w_mem[2344] = 222;
razn_w_mem[2345] = 222;
razn_w_mem[2346] = 222;
razn_w_mem[2347] = 222;
razn_w_mem[2348] = 222;
razn_w_mem[2349] = 222;
razn_w_mem[2350] = 222;
razn_w_mem[2351] = 222;
razn_w_mem[2352] = 222;
razn_w_mem[2353] = 222;
razn_w_mem[2354] = 222;
razn_w_mem[2355] = 222;
razn_w_mem[2356] = 222;
razn_w_mem[2357] = 222;
razn_w_mem[2358] = 222;
razn_w_mem[2359] = 222;
razn_w_mem[2360] = 222;
razn_w_mem[2361] = 222;
razn_w_mem[2362] = 222;
razn_w_mem[2363] = 222;
razn_w_mem[2364] = 222;
razn_w_mem[2365] = 222;
razn_w_mem[2366] = 222;
razn_w_mem[2367] = 222;
razn_w_mem[2368] = 222;
razn_w_mem[2369] = 222;
razn_w_mem[2370] = 222;
razn_w_mem[2371] = 222;
razn_w_mem[2372] = 222;
razn_w_mem[2373] = 222;
razn_w_mem[2374] = 222;
razn_w_mem[2375] = 222;
razn_w_mem[2376] = 222;
razn_w_mem[2377] = 222;
razn_w_mem[2378] = 222;
razn_w_mem[2379] = 222;
razn_w_mem[2380] = 222;
razn_w_mem[2381] = 222;
razn_w_mem[2382] = 222;
razn_w_mem[2383] = 222;
razn_w_mem[2384] = 222;
razn_w_mem[2385] = 222;
razn_w_mem[2386] = 222;
razn_w_mem[2387] = 222;
razn_w_mem[2388] = 222;
razn_w_mem[2389] = 222;
razn_w_mem[2390] = 222;
razn_w_mem[2391] = 222;
razn_w_mem[2392] = 222;
razn_w_mem[2393] = 222;
razn_w_mem[2394] = 222;
razn_w_mem[2395] = 222;
razn_w_mem[2396] = 222;
razn_w_mem[2397] = 222;
razn_w_mem[2398] = 222;
razn_w_mem[2399] = 222;
razn_w_mem[2400] = 222;
razn_w_mem[2401] = 222;
razn_w_mem[2402] = 222;
razn_w_mem[2403] = 222;
razn_w_mem[2404] = 222;
razn_w_mem[2405] = 222;
razn_w_mem[2406] = 222;
razn_w_mem[2407] = 222;
razn_w_mem[2408] = 222;
razn_w_mem[2409] = 222;
razn_w_mem[2410] = 222;
razn_w_mem[2411] = 222;
razn_w_mem[2412] = 222;
razn_w_mem[2413] = 222;
razn_w_mem[2414] = 222;
razn_w_mem[2415] = 222;
razn_w_mem[2416] = 222;
razn_w_mem[2417] = 222;
razn_w_mem[2418] = 222;
razn_w_mem[2419] = 222;
razn_w_mem[2420] = 222;
razn_w_mem[2421] = 222;
razn_w_mem[2422] = 222;
razn_w_mem[2423] = 222;
razn_w_mem[2424] = 222;
razn_w_mem[2425] = 222;
razn_w_mem[2426] = 222;
razn_w_mem[2427] = 222;
razn_w_mem[2428] = 222;
razn_w_mem[2429] = 222;
razn_w_mem[2430] = 222;
razn_w_mem[2431] = 222;
razn_w_mem[2432] = 192;
razn_w_mem[2433] = 192;
razn_w_mem[2434] = 192;
razn_w_mem[2435] = 192;
razn_w_mem[2436] = 192;
razn_w_mem[2437] = 192;
razn_w_mem[2438] = 192;
razn_w_mem[2439] = 192;
razn_w_mem[2440] = 192;
razn_w_mem[2441] = 192;
razn_w_mem[2442] = 192;
razn_w_mem[2443] = 192;
razn_w_mem[2444] = 192;
razn_w_mem[2445] = 192;
razn_w_mem[2446] = 192;
razn_w_mem[2447] = 192;
razn_w_mem[2448] = 192;
razn_w_mem[2449] = 192;
razn_w_mem[2450] = 192;
razn_w_mem[2451] = 192;
razn_w_mem[2452] = 192;
razn_w_mem[2453] = 192;
razn_w_mem[2454] = 192;
razn_w_mem[2455] = 192;
razn_w_mem[2456] = 192;
razn_w_mem[2457] = 192;
razn_w_mem[2458] = 192;
razn_w_mem[2459] = 192;
razn_w_mem[2460] = 192;
razn_w_mem[2461] = 192;
razn_w_mem[2462] = 192;
razn_w_mem[2463] = 192;
razn_w_mem[2464] = 192;
razn_w_mem[2465] = 192;
razn_w_mem[2466] = 192;
razn_w_mem[2467] = 192;
razn_w_mem[2468] = 192;
razn_w_mem[2469] = 192;
razn_w_mem[2470] = 192;
razn_w_mem[2471] = 192;
razn_w_mem[2472] = 192;
razn_w_mem[2473] = 192;
razn_w_mem[2474] = 192;
razn_w_mem[2475] = 192;
razn_w_mem[2476] = 192;
razn_w_mem[2477] = 192;
razn_w_mem[2478] = 192;
razn_w_mem[2479] = 192;
razn_w_mem[2480] = 192;
razn_w_mem[2481] = 192;
razn_w_mem[2482] = 192;
razn_w_mem[2483] = 192;
razn_w_mem[2484] = 192;
razn_w_mem[2485] = 192;
razn_w_mem[2486] = 192;
razn_w_mem[2487] = 192;
razn_w_mem[2488] = 192;
razn_w_mem[2489] = 192;
razn_w_mem[2490] = 192;
razn_w_mem[2491] = 192;
razn_w_mem[2492] = 192;
razn_w_mem[2493] = 192;
razn_w_mem[2494] = 192;
razn_w_mem[2495] = 192;
razn_w_mem[2496] = 192;
razn_w_mem[2497] = 192;
razn_w_mem[2498] = 192;
razn_w_mem[2499] = 192;
razn_w_mem[2500] = 192;
razn_w_mem[2501] = 192;
razn_w_mem[2502] = 192;
razn_w_mem[2503] = 192;
razn_w_mem[2504] = 192;
razn_w_mem[2505] = 192;
razn_w_mem[2506] = 192;
razn_w_mem[2507] = 192;
razn_w_mem[2508] = 192;
razn_w_mem[2509] = 192;
razn_w_mem[2510] = 192;
razn_w_mem[2511] = 192;
razn_w_mem[2512] = 192;
razn_w_mem[2513] = 192;
razn_w_mem[2514] = 192;
razn_w_mem[2515] = 192;
razn_w_mem[2516] = 192;
razn_w_mem[2517] = 192;
razn_w_mem[2518] = 192;
razn_w_mem[2519] = 192;
razn_w_mem[2520] = 192;
razn_w_mem[2521] = 192;
razn_w_mem[2522] = 192;
razn_w_mem[2523] = 192;
razn_w_mem[2524] = 192;
razn_w_mem[2525] = 192;
razn_w_mem[2526] = 192;
razn_w_mem[2527] = 192;
razn_w_mem[2528] = 192;
razn_w_mem[2529] = 192;
razn_w_mem[2530] = 192;
razn_w_mem[2531] = 192;
razn_w_mem[2532] = 192;
razn_w_mem[2533] = 192;
razn_w_mem[2534] = 192;
razn_w_mem[2535] = 192;
razn_w_mem[2536] = 192;
razn_w_mem[2537] = 192;
razn_w_mem[2538] = 192;
razn_w_mem[2539] = 192;
razn_w_mem[2540] = 192;
razn_w_mem[2541] = 192;
razn_w_mem[2542] = 192;
razn_w_mem[2543] = 192;
razn_w_mem[2544] = 192;
razn_w_mem[2545] = 192;
razn_w_mem[2546] = 192;
razn_w_mem[2547] = 192;
razn_w_mem[2548] = 192;
razn_w_mem[2549] = 192;
razn_w_mem[2550] = 192;
razn_w_mem[2551] = 192;
razn_w_mem[2552] = 192;
razn_w_mem[2553] = 192;
razn_w_mem[2554] = 192;
razn_w_mem[2555] = 192;
razn_w_mem[2556] = 192;
razn_w_mem[2557] = 192;
razn_w_mem[2558] = 192;
razn_w_mem[2559] = 192;
razn_w_mem[2560] = 162;
razn_w_mem[2561] = 162;
razn_w_mem[2562] = 162;
razn_w_mem[2563] = 162;
razn_w_mem[2564] = 162;
razn_w_mem[2565] = 162;
razn_w_mem[2566] = 162;
razn_w_mem[2567] = 162;
razn_w_mem[2568] = 162;
razn_w_mem[2569] = 162;
razn_w_mem[2570] = 162;
razn_w_mem[2571] = 162;
razn_w_mem[2572] = 162;
razn_w_mem[2573] = 162;
razn_w_mem[2574] = 162;
razn_w_mem[2575] = 162;
razn_w_mem[2576] = 162;
razn_w_mem[2577] = 162;
razn_w_mem[2578] = 162;
razn_w_mem[2579] = 162;
razn_w_mem[2580] = 162;
razn_w_mem[2581] = 162;
razn_w_mem[2582] = 162;
razn_w_mem[2583] = 162;
razn_w_mem[2584] = 162;
razn_w_mem[2585] = 162;
razn_w_mem[2586] = 162;
razn_w_mem[2587] = 162;
razn_w_mem[2588] = 162;
razn_w_mem[2589] = 162;
razn_w_mem[2590] = 162;
razn_w_mem[2591] = 162;
razn_w_mem[2592] = 162;
razn_w_mem[2593] = 162;
razn_w_mem[2594] = 162;
razn_w_mem[2595] = 162;
razn_w_mem[2596] = 162;
razn_w_mem[2597] = 162;
razn_w_mem[2598] = 162;
razn_w_mem[2599] = 162;
razn_w_mem[2600] = 162;
razn_w_mem[2601] = 162;
razn_w_mem[2602] = 162;
razn_w_mem[2603] = 162;
razn_w_mem[2604] = 162;
razn_w_mem[2605] = 162;
razn_w_mem[2606] = 162;
razn_w_mem[2607] = 162;
razn_w_mem[2608] = 162;
razn_w_mem[2609] = 162;
razn_w_mem[2610] = 162;
razn_w_mem[2611] = 162;
razn_w_mem[2612] = 162;
razn_w_mem[2613] = 162;
razn_w_mem[2614] = 162;
razn_w_mem[2615] = 162;
razn_w_mem[2616] = 162;
razn_w_mem[2617] = 162;
razn_w_mem[2618] = 162;
razn_w_mem[2619] = 162;
razn_w_mem[2620] = 162;
razn_w_mem[2621] = 162;
razn_w_mem[2622] = 162;
razn_w_mem[2623] = 162;
razn_w_mem[2624] = 162;
razn_w_mem[2625] = 162;
razn_w_mem[2626] = 162;
razn_w_mem[2627] = 162;
razn_w_mem[2628] = 162;
razn_w_mem[2629] = 162;
razn_w_mem[2630] = 162;
razn_w_mem[2631] = 162;
razn_w_mem[2632] = 162;
razn_w_mem[2633] = 162;
razn_w_mem[2634] = 162;
razn_w_mem[2635] = 162;
razn_w_mem[2636] = 162;
razn_w_mem[2637] = 162;
razn_w_mem[2638] = 162;
razn_w_mem[2639] = 162;
razn_w_mem[2640] = 162;
razn_w_mem[2641] = 162;
razn_w_mem[2642] = 162;
razn_w_mem[2643] = 162;
razn_w_mem[2644] = 162;
razn_w_mem[2645] = 162;
razn_w_mem[2646] = 162;
razn_w_mem[2647] = 162;
razn_w_mem[2648] = 162;
razn_w_mem[2649] = 162;
razn_w_mem[2650] = 162;
razn_w_mem[2651] = 162;
razn_w_mem[2652] = 162;
razn_w_mem[2653] = 162;
razn_w_mem[2654] = 162;
razn_w_mem[2655] = 162;
razn_w_mem[2656] = 162;
razn_w_mem[2657] = 162;
razn_w_mem[2658] = 162;
razn_w_mem[2659] = 162;
razn_w_mem[2660] = 162;
razn_w_mem[2661] = 162;
razn_w_mem[2662] = 162;
razn_w_mem[2663] = 162;
razn_w_mem[2664] = 162;
razn_w_mem[2665] = 162;
razn_w_mem[2666] = 162;
razn_w_mem[2667] = 162;
razn_w_mem[2668] = 162;
razn_w_mem[2669] = 162;
razn_w_mem[2670] = 162;
razn_w_mem[2671] = 162;
razn_w_mem[2672] = 162;
razn_w_mem[2673] = 162;
razn_w_mem[2674] = 162;
razn_w_mem[2675] = 162;
razn_w_mem[2676] = 162;
razn_w_mem[2677] = 162;
razn_w_mem[2678] = 162;
razn_w_mem[2679] = 162;
razn_w_mem[2680] = 162;
razn_w_mem[2681] = 162;
razn_w_mem[2682] = 162;
razn_w_mem[2683] = 162;
razn_w_mem[2684] = 162;
razn_w_mem[2685] = 162;
razn_w_mem[2686] = 162;
razn_w_mem[2687] = 162;
razn_w_mem[2688] = 132;
razn_w_mem[2689] = 132;
razn_w_mem[2690] = 132;
razn_w_mem[2691] = 132;
razn_w_mem[2692] = 132;
razn_w_mem[2693] = 132;
razn_w_mem[2694] = 132;
razn_w_mem[2695] = 132;
razn_w_mem[2696] = 132;
razn_w_mem[2697] = 132;
razn_w_mem[2698] = 132;
razn_w_mem[2699] = 132;
razn_w_mem[2700] = 132;
razn_w_mem[2701] = 132;
razn_w_mem[2702] = 132;
razn_w_mem[2703] = 132;
razn_w_mem[2704] = 132;
razn_w_mem[2705] = 132;
razn_w_mem[2706] = 132;
razn_w_mem[2707] = 132;
razn_w_mem[2708] = 132;
razn_w_mem[2709] = 132;
razn_w_mem[2710] = 132;
razn_w_mem[2711] = 132;
razn_w_mem[2712] = 132;
razn_w_mem[2713] = 132;
razn_w_mem[2714] = 132;
razn_w_mem[2715] = 132;
razn_w_mem[2716] = 132;
razn_w_mem[2717] = 132;
razn_w_mem[2718] = 132;
razn_w_mem[2719] = 132;
razn_w_mem[2720] = 132;
razn_w_mem[2721] = 132;
razn_w_mem[2722] = 132;
razn_w_mem[2723] = 132;
razn_w_mem[2724] = 132;
razn_w_mem[2725] = 132;
razn_w_mem[2726] = 132;
razn_w_mem[2727] = 132;
razn_w_mem[2728] = 132;
razn_w_mem[2729] = 132;
razn_w_mem[2730] = 132;
razn_w_mem[2731] = 132;
razn_w_mem[2732] = 132;
razn_w_mem[2733] = 132;
razn_w_mem[2734] = 132;
razn_w_mem[2735] = 132;
razn_w_mem[2736] = 132;
razn_w_mem[2737] = 132;
razn_w_mem[2738] = 132;
razn_w_mem[2739] = 132;
razn_w_mem[2740] = 132;
razn_w_mem[2741] = 132;
razn_w_mem[2742] = 132;
razn_w_mem[2743] = 132;
razn_w_mem[2744] = 132;
razn_w_mem[2745] = 132;
razn_w_mem[2746] = 132;
razn_w_mem[2747] = 132;
razn_w_mem[2748] = 132;
razn_w_mem[2749] = 132;
razn_w_mem[2750] = 132;
razn_w_mem[2751] = 132;
razn_w_mem[2752] = 132;
razn_w_mem[2753] = 132;
razn_w_mem[2754] = 132;
razn_w_mem[2755] = 132;
razn_w_mem[2756] = 132;
razn_w_mem[2757] = 132;
razn_w_mem[2758] = 132;
razn_w_mem[2759] = 132;
razn_w_mem[2760] = 132;
razn_w_mem[2761] = 132;
razn_w_mem[2762] = 132;
razn_w_mem[2763] = 132;
razn_w_mem[2764] = 132;
razn_w_mem[2765] = 132;
razn_w_mem[2766] = 132;
razn_w_mem[2767] = 132;
razn_w_mem[2768] = 132;
razn_w_mem[2769] = 132;
razn_w_mem[2770] = 132;
razn_w_mem[2771] = 132;
razn_w_mem[2772] = 132;
razn_w_mem[2773] = 132;
razn_w_mem[2774] = 132;
razn_w_mem[2775] = 132;
razn_w_mem[2776] = 132;
razn_w_mem[2777] = 132;
razn_w_mem[2778] = 132;
razn_w_mem[2779] = 132;
razn_w_mem[2780] = 132;
razn_w_mem[2781] = 132;
razn_w_mem[2782] = 132;
razn_w_mem[2783] = 132;
razn_w_mem[2784] = 132;
razn_w_mem[2785] = 132;
razn_w_mem[2786] = 132;
razn_w_mem[2787] = 132;
razn_w_mem[2788] = 132;
razn_w_mem[2789] = 132;
razn_w_mem[2790] = 132;
razn_w_mem[2791] = 132;
razn_w_mem[2792] = 132;
razn_w_mem[2793] = 132;
razn_w_mem[2794] = 132;
razn_w_mem[2795] = 132;
razn_w_mem[2796] = 132;
razn_w_mem[2797] = 132;
razn_w_mem[2798] = 132;
razn_w_mem[2799] = 132;
razn_w_mem[2800] = 132;
razn_w_mem[2801] = 132;
razn_w_mem[2802] = 132;
razn_w_mem[2803] = 132;
razn_w_mem[2804] = 132;
razn_w_mem[2805] = 132;
razn_w_mem[2806] = 132;
razn_w_mem[2807] = 132;
razn_w_mem[2808] = 132;
razn_w_mem[2809] = 132;
razn_w_mem[2810] = 132;
razn_w_mem[2811] = 132;
razn_w_mem[2812] = 132;
razn_w_mem[2813] = 132;
razn_w_mem[2814] = 132;
razn_w_mem[2815] = 132;
razn_w_mem[2816] = 102;
razn_w_mem[2817] = 102;
razn_w_mem[2818] = 102;
razn_w_mem[2819] = 102;
razn_w_mem[2820] = 102;
razn_w_mem[2821] = 102;
razn_w_mem[2822] = 102;
razn_w_mem[2823] = 102;
razn_w_mem[2824] = 102;
razn_w_mem[2825] = 102;
razn_w_mem[2826] = 102;
razn_w_mem[2827] = 102;
razn_w_mem[2828] = 102;
razn_w_mem[2829] = 102;
razn_w_mem[2830] = 102;
razn_w_mem[2831] = 102;
razn_w_mem[2832] = 102;
razn_w_mem[2833] = 102;
razn_w_mem[2834] = 102;
razn_w_mem[2835] = 102;
razn_w_mem[2836] = 102;
razn_w_mem[2837] = 102;
razn_w_mem[2838] = 102;
razn_w_mem[2839] = 102;
razn_w_mem[2840] = 102;
razn_w_mem[2841] = 102;
razn_w_mem[2842] = 102;
razn_w_mem[2843] = 102;
razn_w_mem[2844] = 102;
razn_w_mem[2845] = 102;
razn_w_mem[2846] = 102;
razn_w_mem[2847] = 102;
razn_w_mem[2848] = 102;
razn_w_mem[2849] = 102;
razn_w_mem[2850] = 102;
razn_w_mem[2851] = 102;
razn_w_mem[2852] = 102;
razn_w_mem[2853] = 102;
razn_w_mem[2854] = 102;
razn_w_mem[2855] = 102;
razn_w_mem[2856] = 102;
razn_w_mem[2857] = 102;
razn_w_mem[2858] = 102;
razn_w_mem[2859] = 102;
razn_w_mem[2860] = 102;
razn_w_mem[2861] = 102;
razn_w_mem[2862] = 102;
razn_w_mem[2863] = 102;
razn_w_mem[2864] = 102;
razn_w_mem[2865] = 102;
razn_w_mem[2866] = 102;
razn_w_mem[2867] = 102;
razn_w_mem[2868] = 102;
razn_w_mem[2869] = 102;
razn_w_mem[2870] = 102;
razn_w_mem[2871] = 102;
razn_w_mem[2872] = 102;
razn_w_mem[2873] = 102;
razn_w_mem[2874] = 102;
razn_w_mem[2875] = 102;
razn_w_mem[2876] = 102;
razn_w_mem[2877] = 102;
razn_w_mem[2878] = 102;
razn_w_mem[2879] = 102;
razn_w_mem[2880] = 102;
razn_w_mem[2881] = 102;
razn_w_mem[2882] = 102;
razn_w_mem[2883] = 102;
razn_w_mem[2884] = 102;
razn_w_mem[2885] = 102;
razn_w_mem[2886] = 102;
razn_w_mem[2887] = 102;
razn_w_mem[2888] = 102;
razn_w_mem[2889] = 102;
razn_w_mem[2890] = 102;
razn_w_mem[2891] = 102;
razn_w_mem[2892] = 102;
razn_w_mem[2893] = 102;
razn_w_mem[2894] = 102;
razn_w_mem[2895] = 102;
razn_w_mem[2896] = 102;
razn_w_mem[2897] = 102;
razn_w_mem[2898] = 102;
razn_w_mem[2899] = 102;
razn_w_mem[2900] = 102;
razn_w_mem[2901] = 102;
razn_w_mem[2902] = 102;
razn_w_mem[2903] = 102;
razn_w_mem[2904] = 102;
razn_w_mem[2905] = 102;
razn_w_mem[2906] = 102;
razn_w_mem[2907] = 102;
razn_w_mem[2908] = 102;
razn_w_mem[2909] = 102;
razn_w_mem[2910] = 102;
razn_w_mem[2911] = 102;
razn_w_mem[2912] = 102;
razn_w_mem[2913] = 102;
razn_w_mem[2914] = 102;
razn_w_mem[2915] = 102;
razn_w_mem[2916] = 102;
razn_w_mem[2917] = 102;
razn_w_mem[2918] = 102;
razn_w_mem[2919] = 102;
razn_w_mem[2920] = 102;
razn_w_mem[2921] = 102;
razn_w_mem[2922] = 102;
razn_w_mem[2923] = 102;
razn_w_mem[2924] = 102;
razn_w_mem[2925] = 102;
razn_w_mem[2926] = 102;
razn_w_mem[2927] = 102;
razn_w_mem[2928] = 102;
razn_w_mem[2929] = 102;
razn_w_mem[2930] = 102;
razn_w_mem[2931] = 102;
razn_w_mem[2932] = 102;
razn_w_mem[2933] = 102;
razn_w_mem[2934] = 102;
razn_w_mem[2935] = 102;
razn_w_mem[2936] = 102;
razn_w_mem[2937] = 102;
razn_w_mem[2938] = 102;
razn_w_mem[2939] = 102;
razn_w_mem[2940] = 102;
razn_w_mem[2941] = 102;
razn_w_mem[2942] = 102;
razn_w_mem[2943] = 102;
razn_w_mem[2944] = 72;
razn_w_mem[2945] = 72;
razn_w_mem[2946] = 72;
razn_w_mem[2947] = 72;
razn_w_mem[2948] = 72;
razn_w_mem[2949] = 72;
razn_w_mem[2950] = 72;
razn_w_mem[2951] = 72;
razn_w_mem[2952] = 72;
razn_w_mem[2953] = 72;
razn_w_mem[2954] = 72;
razn_w_mem[2955] = 72;
razn_w_mem[2956] = 72;
razn_w_mem[2957] = 72;
razn_w_mem[2958] = 72;
razn_w_mem[2959] = 72;
razn_w_mem[2960] = 72;
razn_w_mem[2961] = 72;
razn_w_mem[2962] = 72;
razn_w_mem[2963] = 72;
razn_w_mem[2964] = 72;
razn_w_mem[2965] = 72;
razn_w_mem[2966] = 72;
razn_w_mem[2967] = 72;
razn_w_mem[2968] = 72;
razn_w_mem[2969] = 72;
razn_w_mem[2970] = 72;
razn_w_mem[2971] = 72;
razn_w_mem[2972] = 72;
razn_w_mem[2973] = 72;
razn_w_mem[2974] = 72;
razn_w_mem[2975] = 72;
razn_w_mem[2976] = 72;
razn_w_mem[2977] = 72;
razn_w_mem[2978] = 72;
razn_w_mem[2979] = 72;
razn_w_mem[2980] = 72;
razn_w_mem[2981] = 72;
razn_w_mem[2982] = 72;
razn_w_mem[2983] = 72;
razn_w_mem[2984] = 72;
razn_w_mem[2985] = 72;
razn_w_mem[2986] = 72;
razn_w_mem[2987] = 72;
razn_w_mem[2988] = 72;
razn_w_mem[2989] = 72;
razn_w_mem[2990] = 72;
razn_w_mem[2991] = 72;
razn_w_mem[2992] = 72;
razn_w_mem[2993] = 72;
razn_w_mem[2994] = 72;
razn_w_mem[2995] = 72;
razn_w_mem[2996] = 72;
razn_w_mem[2997] = 72;
razn_w_mem[2998] = 72;
razn_w_mem[2999] = 72;
razn_w_mem[3000] = 72;
razn_w_mem[3001] = 72;
razn_w_mem[3002] = 72;
razn_w_mem[3003] = 72;
razn_w_mem[3004] = 72;
razn_w_mem[3005] = 72;
razn_w_mem[3006] = 72;
razn_w_mem[3007] = 72;
razn_w_mem[3008] = 72;
razn_w_mem[3009] = 72;
razn_w_mem[3010] = 72;
razn_w_mem[3011] = 72;
razn_w_mem[3012] = 72;
razn_w_mem[3013] = 72;
razn_w_mem[3014] = 72;
razn_w_mem[3015] = 72;
razn_w_mem[3016] = 72;
razn_w_mem[3017] = 72;
razn_w_mem[3018] = 72;
razn_w_mem[3019] = 72;
razn_w_mem[3020] = 72;
razn_w_mem[3021] = 72;
razn_w_mem[3022] = 72;
razn_w_mem[3023] = 72;
razn_w_mem[3024] = 72;
razn_w_mem[3025] = 72;
razn_w_mem[3026] = 72;
razn_w_mem[3027] = 72;
razn_w_mem[3028] = 72;
razn_w_mem[3029] = 72;
razn_w_mem[3030] = 72;
razn_w_mem[3031] = 72;
razn_w_mem[3032] = 72;
razn_w_mem[3033] = 72;
razn_w_mem[3034] = 72;
razn_w_mem[3035] = 72;
razn_w_mem[3036] = 72;
razn_w_mem[3037] = 72;
razn_w_mem[3038] = 72;
razn_w_mem[3039] = 72;
razn_w_mem[3040] = 72;
razn_w_mem[3041] = 72;
razn_w_mem[3042] = 72;
razn_w_mem[3043] = 72;
razn_w_mem[3044] = 72;
razn_w_mem[3045] = 72;
razn_w_mem[3046] = 72;
razn_w_mem[3047] = 72;
razn_w_mem[3048] = 72;
razn_w_mem[3049] = 72;
razn_w_mem[3050] = 72;
razn_w_mem[3051] = 72;
razn_w_mem[3052] = 72;
razn_w_mem[3053] = 72;
razn_w_mem[3054] = 72;
razn_w_mem[3055] = 72;
razn_w_mem[3056] = 72;
razn_w_mem[3057] = 72;
razn_w_mem[3058] = 72;
razn_w_mem[3059] = 72;
razn_w_mem[3060] = 72;
razn_w_mem[3061] = 72;
razn_w_mem[3062] = 72;
razn_w_mem[3063] = 72;
razn_w_mem[3064] = 72;
razn_w_mem[3065] = 72;
razn_w_mem[3066] = 72;
razn_w_mem[3067] = 72;
razn_w_mem[3068] = 72;
razn_w_mem[3069] = 72;
razn_w_mem[3070] = 72;
razn_w_mem[3071] = 72;
razn_w_mem[3072] = 42;
razn_w_mem[3073] = 42;
razn_w_mem[3074] = 42;
razn_w_mem[3075] = 42;
razn_w_mem[3076] = 42;
razn_w_mem[3077] = 42;
razn_w_mem[3078] = 42;
razn_w_mem[3079] = 42;
razn_w_mem[3080] = 42;
razn_w_mem[3081] = 42;
razn_w_mem[3082] = 42;
razn_w_mem[3083] = 42;
razn_w_mem[3084] = 42;
razn_w_mem[3085] = 42;
razn_w_mem[3086] = 42;
razn_w_mem[3087] = 42;
razn_w_mem[3088] = 42;
razn_w_mem[3089] = 42;
razn_w_mem[3090] = 42;
razn_w_mem[3091] = 42;
razn_w_mem[3092] = 42;
razn_w_mem[3093] = 42;
razn_w_mem[3094] = 42;
razn_w_mem[3095] = 42;
razn_w_mem[3096] = 42;
razn_w_mem[3097] = 42;
razn_w_mem[3098] = 42;
razn_w_mem[3099] = 42;
razn_w_mem[3100] = 42;
razn_w_mem[3101] = 42;
razn_w_mem[3102] = 42;
razn_w_mem[3103] = 42;
razn_w_mem[3104] = 42;
razn_w_mem[3105] = 42;
razn_w_mem[3106] = 42;
razn_w_mem[3107] = 42;
razn_w_mem[3108] = 42;
razn_w_mem[3109] = 42;
razn_w_mem[3110] = 42;
razn_w_mem[3111] = 42;
razn_w_mem[3112] = 42;
razn_w_mem[3113] = 42;
razn_w_mem[3114] = 42;
razn_w_mem[3115] = 42;
razn_w_mem[3116] = 42;
razn_w_mem[3117] = 42;
razn_w_mem[3118] = 42;
razn_w_mem[3119] = 42;
razn_w_mem[3120] = 42;
razn_w_mem[3121] = 42;
razn_w_mem[3122] = 42;
razn_w_mem[3123] = 42;
razn_w_mem[3124] = 42;
razn_w_mem[3125] = 42;
razn_w_mem[3126] = 42;
razn_w_mem[3127] = 42;
razn_w_mem[3128] = 42;
razn_w_mem[3129] = 42;
razn_w_mem[3130] = 42;
razn_w_mem[3131] = 42;
razn_w_mem[3132] = 42;
razn_w_mem[3133] = 42;
razn_w_mem[3134] = 42;
razn_w_mem[3135] = 42;
razn_w_mem[3136] = 42;
razn_w_mem[3137] = 42;
razn_w_mem[3138] = 42;
razn_w_mem[3139] = 42;
razn_w_mem[3140] = 42;
razn_w_mem[3141] = 42;
razn_w_mem[3142] = 42;
razn_w_mem[3143] = 42;
razn_w_mem[3144] = 42;
razn_w_mem[3145] = 42;
razn_w_mem[3146] = 42;
razn_w_mem[3147] = 42;
razn_w_mem[3148] = 42;
razn_w_mem[3149] = 42;
razn_w_mem[3150] = 42;
razn_w_mem[3151] = 42;
razn_w_mem[3152] = 42;
razn_w_mem[3153] = 42;
razn_w_mem[3154] = 42;
razn_w_mem[3155] = 42;
razn_w_mem[3156] = 42;
razn_w_mem[3157] = 42;
razn_w_mem[3158] = 42;
razn_w_mem[3159] = 42;
razn_w_mem[3160] = 42;
razn_w_mem[3161] = 42;
razn_w_mem[3162] = 42;
razn_w_mem[3163] = 42;
razn_w_mem[3164] = 42;
razn_w_mem[3165] = 42;
razn_w_mem[3166] = 42;
razn_w_mem[3167] = 42;
razn_w_mem[3168] = 42;
razn_w_mem[3169] = 42;
razn_w_mem[3170] = 42;
razn_w_mem[3171] = 42;
razn_w_mem[3172] = 42;
razn_w_mem[3173] = 42;
razn_w_mem[3174] = 42;
razn_w_mem[3175] = 42;
razn_w_mem[3176] = 42;
razn_w_mem[3177] = 42;
razn_w_mem[3178] = 42;
razn_w_mem[3179] = 42;
razn_w_mem[3180] = 42;
razn_w_mem[3181] = 42;
razn_w_mem[3182] = 42;
razn_w_mem[3183] = 42;
razn_w_mem[3184] = 42;
razn_w_mem[3185] = 42;
razn_w_mem[3186] = 42;
razn_w_mem[3187] = 42;
razn_w_mem[3188] = 42;
razn_w_mem[3189] = 42;
razn_w_mem[3190] = 42;
razn_w_mem[3191] = 42;
razn_w_mem[3192] = 42;
razn_w_mem[3193] = 42;
razn_w_mem[3194] = 42;
razn_w_mem[3195] = 42;
razn_w_mem[3196] = 42;
razn_w_mem[3197] = 42;
razn_w_mem[3198] = 42;
razn_w_mem[3199] = 42;
razn_w_mem[3200] = 12;
razn_w_mem[3201] = 12;
razn_w_mem[3202] = 12;
razn_w_mem[3203] = 12;
razn_w_mem[3204] = 12;
razn_w_mem[3205] = 12;
razn_w_mem[3206] = 12;
razn_w_mem[3207] = 12;
razn_w_mem[3208] = 12;
razn_w_mem[3209] = 12;
razn_w_mem[3210] = 12;
razn_w_mem[3211] = 12;
razn_w_mem[3212] = 12;
razn_w_mem[3213] = 12;
razn_w_mem[3214] = 12;
razn_w_mem[3215] = 12;
razn_w_mem[3216] = 12;
razn_w_mem[3217] = 12;
razn_w_mem[3218] = 12;
razn_w_mem[3219] = 12;
razn_w_mem[3220] = 12;
razn_w_mem[3221] = 12;
razn_w_mem[3222] = 12;
razn_w_mem[3223] = 12;
razn_w_mem[3224] = 12;
razn_w_mem[3225] = 12;
razn_w_mem[3226] = 12;
razn_w_mem[3227] = 12;
razn_w_mem[3228] = 12;
razn_w_mem[3229] = 12;
razn_w_mem[3230] = 12;
razn_w_mem[3231] = 12;
razn_w_mem[3232] = 12;
razn_w_mem[3233] = 12;
razn_w_mem[3234] = 12;
razn_w_mem[3235] = 12;
razn_w_mem[3236] = 12;
razn_w_mem[3237] = 12;
razn_w_mem[3238] = 12;
razn_w_mem[3239] = 12;
razn_w_mem[3240] = 12;
razn_w_mem[3241] = 12;
razn_w_mem[3242] = 12;
razn_w_mem[3243] = 12;
razn_w_mem[3244] = 12;
razn_w_mem[3245] = 12;
razn_w_mem[3246] = 12;
razn_w_mem[3247] = 12;
razn_w_mem[3248] = 12;
razn_w_mem[3249] = 12;
razn_w_mem[3250] = 12;
razn_w_mem[3251] = 12;
razn_w_mem[3252] = 12;
razn_w_mem[3253] = 12;
razn_w_mem[3254] = 12;
razn_w_mem[3255] = 12;
razn_w_mem[3256] = 12;
razn_w_mem[3257] = 12;
razn_w_mem[3258] = 12;
razn_w_mem[3259] = 12;
razn_w_mem[3260] = 12;
razn_w_mem[3261] = 12;
razn_w_mem[3262] = 12;
razn_w_mem[3263] = 12;
razn_w_mem[3264] = 12;
razn_w_mem[3265] = 12;
razn_w_mem[3266] = 12;
razn_w_mem[3267] = 12;
razn_w_mem[3268] = 12;
razn_w_mem[3269] = 12;
razn_w_mem[3270] = 12;
razn_w_mem[3271] = 12;
razn_w_mem[3272] = 12;
razn_w_mem[3273] = 12;
razn_w_mem[3274] = 12;
razn_w_mem[3275] = 12;
razn_w_mem[3276] = 12;
razn_w_mem[3277] = 12;
razn_w_mem[3278] = 12;
razn_w_mem[3279] = 12;
razn_w_mem[3280] = 12;
razn_w_mem[3281] = 12;
razn_w_mem[3282] = 12;
razn_w_mem[3283] = 12;
razn_w_mem[3284] = 12;
razn_w_mem[3285] = 12;
razn_w_mem[3286] = 12;
razn_w_mem[3287] = 12;
razn_w_mem[3288] = 12;
razn_w_mem[3289] = 12;
razn_w_mem[3290] = 12;
razn_w_mem[3291] = 12;
razn_w_mem[3292] = 12;
razn_w_mem[3293] = 12;
razn_w_mem[3294] = 12;
razn_w_mem[3295] = 12;
razn_w_mem[3296] = 12;
razn_w_mem[3297] = 12;
razn_w_mem[3298] = 12;
razn_w_mem[3299] = 12;
razn_w_mem[3300] = 12;
razn_w_mem[3301] = 12;
razn_w_mem[3302] = 12;
razn_w_mem[3303] = 12;
razn_w_mem[3304] = 12;
razn_w_mem[3305] = 12;
razn_w_mem[3306] = 12;
razn_w_mem[3307] = 12;
razn_w_mem[3308] = 12;
razn_w_mem[3309] = 12;
razn_w_mem[3310] = 12;
razn_w_mem[3311] = 12;
razn_w_mem[3312] = 12;
razn_w_mem[3313] = 12;
razn_w_mem[3314] = 12;
razn_w_mem[3315] = 12;
razn_w_mem[3316] = 12;
razn_w_mem[3317] = 12;
razn_w_mem[3318] = 12;
razn_w_mem[3319] = 12;
razn_w_mem[3320] = 12;
razn_w_mem[3321] = 12;
razn_w_mem[3322] = 12;
razn_w_mem[3323] = 12;
razn_w_mem[3324] = 12;
razn_w_mem[3325] = 12;
razn_w_mem[3326] = 12;
razn_w_mem[3327] = 12;
razn_w_mem[3328] = 236;
razn_w_mem[3329] = 236;
razn_w_mem[3330] = 236;
razn_w_mem[3331] = 236;
razn_w_mem[3332] = 236;
razn_w_mem[3333] = 236;
razn_w_mem[3334] = 236;
razn_w_mem[3335] = 236;
razn_w_mem[3336] = 236;
razn_w_mem[3337] = 236;
razn_w_mem[3338] = 236;
razn_w_mem[3339] = 236;
razn_w_mem[3340] = 236;
razn_w_mem[3341] = 236;
razn_w_mem[3342] = 236;
razn_w_mem[3343] = 236;
razn_w_mem[3344] = 236;
razn_w_mem[3345] = 236;
razn_w_mem[3346] = 236;
razn_w_mem[3347] = 236;
razn_w_mem[3348] = 236;
razn_w_mem[3349] = 236;
razn_w_mem[3350] = 236;
razn_w_mem[3351] = 236;
razn_w_mem[3352] = 236;
razn_w_mem[3353] = 236;
razn_w_mem[3354] = 236;
razn_w_mem[3355] = 236;
razn_w_mem[3356] = 236;
razn_w_mem[3357] = 236;
razn_w_mem[3358] = 236;
razn_w_mem[3359] = 236;
razn_w_mem[3360] = 236;
razn_w_mem[3361] = 236;
razn_w_mem[3362] = 236;
razn_w_mem[3363] = 236;
razn_w_mem[3364] = 236;
razn_w_mem[3365] = 236;
razn_w_mem[3366] = 236;
razn_w_mem[3367] = 236;
razn_w_mem[3368] = 236;
razn_w_mem[3369] = 236;
razn_w_mem[3370] = 236;
razn_w_mem[3371] = 236;
razn_w_mem[3372] = 236;
razn_w_mem[3373] = 236;
razn_w_mem[3374] = 236;
razn_w_mem[3375] = 236;
razn_w_mem[3376] = 236;
razn_w_mem[3377] = 236;
razn_w_mem[3378] = 236;
razn_w_mem[3379] = 236;
razn_w_mem[3380] = 236;
razn_w_mem[3381] = 236;
razn_w_mem[3382] = 236;
razn_w_mem[3383] = 236;
razn_w_mem[3384] = 236;
razn_w_mem[3385] = 236;
razn_w_mem[3386] = 236;
razn_w_mem[3387] = 236;
razn_w_mem[3388] = 236;
razn_w_mem[3389] = 236;
razn_w_mem[3390] = 236;
razn_w_mem[3391] = 236;
razn_w_mem[3392] = 236;
razn_w_mem[3393] = 236;
razn_w_mem[3394] = 236;
razn_w_mem[3395] = 236;
razn_w_mem[3396] = 236;
razn_w_mem[3397] = 236;
razn_w_mem[3398] = 236;
razn_w_mem[3399] = 236;
razn_w_mem[3400] = 236;
razn_w_mem[3401] = 236;
razn_w_mem[3402] = 236;
razn_w_mem[3403] = 236;
razn_w_mem[3404] = 236;
razn_w_mem[3405] = 236;
razn_w_mem[3406] = 236;
razn_w_mem[3407] = 236;
razn_w_mem[3408] = 236;
razn_w_mem[3409] = 236;
razn_w_mem[3410] = 236;
razn_w_mem[3411] = 236;
razn_w_mem[3412] = 236;
razn_w_mem[3413] = 236;
razn_w_mem[3414] = 236;
razn_w_mem[3415] = 236;
razn_w_mem[3416] = 236;
razn_w_mem[3417] = 236;
razn_w_mem[3418] = 236;
razn_w_mem[3419] = 236;
razn_w_mem[3420] = 236;
razn_w_mem[3421] = 236;
razn_w_mem[3422] = 236;
razn_w_mem[3423] = 236;
razn_w_mem[3424] = 236;
razn_w_mem[3425] = 236;
razn_w_mem[3426] = 236;
razn_w_mem[3427] = 236;
razn_w_mem[3428] = 236;
razn_w_mem[3429] = 236;
razn_w_mem[3430] = 236;
razn_w_mem[3431] = 236;
razn_w_mem[3432] = 236;
razn_w_mem[3433] = 236;
razn_w_mem[3434] = 236;
razn_w_mem[3435] = 236;
razn_w_mem[3436] = 236;
razn_w_mem[3437] = 236;
razn_w_mem[3438] = 236;
razn_w_mem[3439] = 236;
razn_w_mem[3440] = 236;
razn_w_mem[3441] = 236;
razn_w_mem[3442] = 236;
razn_w_mem[3443] = 236;
razn_w_mem[3444] = 236;
razn_w_mem[3445] = 236;
razn_w_mem[3446] = 236;
razn_w_mem[3447] = 236;
razn_w_mem[3448] = 236;
razn_w_mem[3449] = 236;
razn_w_mem[3450] = 236;
razn_w_mem[3451] = 236;
razn_w_mem[3452] = 236;
razn_w_mem[3453] = 236;
razn_w_mem[3454] = 236;
razn_w_mem[3455] = 236;
razn_w_mem[3456] = 206;
razn_w_mem[3457] = 206;
razn_w_mem[3458] = 206;
razn_w_mem[3459] = 206;
razn_w_mem[3460] = 206;
razn_w_mem[3461] = 206;
razn_w_mem[3462] = 206;
razn_w_mem[3463] = 206;
razn_w_mem[3464] = 206;
razn_w_mem[3465] = 206;
razn_w_mem[3466] = 206;
razn_w_mem[3467] = 206;
razn_w_mem[3468] = 206;
razn_w_mem[3469] = 206;
razn_w_mem[3470] = 206;
razn_w_mem[3471] = 206;
razn_w_mem[3472] = 206;
razn_w_mem[3473] = 206;
razn_w_mem[3474] = 206;
razn_w_mem[3475] = 206;
razn_w_mem[3476] = 206;
razn_w_mem[3477] = 206;
razn_w_mem[3478] = 206;
razn_w_mem[3479] = 206;
razn_w_mem[3480] = 206;
razn_w_mem[3481] = 206;
razn_w_mem[3482] = 206;
razn_w_mem[3483] = 206;
razn_w_mem[3484] = 206;
razn_w_mem[3485] = 206;
razn_w_mem[3486] = 206;
razn_w_mem[3487] = 206;
razn_w_mem[3488] = 206;
razn_w_mem[3489] = 206;
razn_w_mem[3490] = 206;
razn_w_mem[3491] = 206;
razn_w_mem[3492] = 206;
razn_w_mem[3493] = 206;
razn_w_mem[3494] = 206;
razn_w_mem[3495] = 206;
razn_w_mem[3496] = 206;
razn_w_mem[3497] = 206;
razn_w_mem[3498] = 206;
razn_w_mem[3499] = 206;
razn_w_mem[3500] = 206;
razn_w_mem[3501] = 206;
razn_w_mem[3502] = 206;
razn_w_mem[3503] = 206;
razn_w_mem[3504] = 206;
razn_w_mem[3505] = 206;
razn_w_mem[3506] = 206;
razn_w_mem[3507] = 206;
razn_w_mem[3508] = 206;
razn_w_mem[3509] = 206;
razn_w_mem[3510] = 206;
razn_w_mem[3511] = 206;
razn_w_mem[3512] = 206;
razn_w_mem[3513] = 206;
razn_w_mem[3514] = 206;
razn_w_mem[3515] = 206;
razn_w_mem[3516] = 206;
razn_w_mem[3517] = 206;
razn_w_mem[3518] = 206;
razn_w_mem[3519] = 206;
razn_w_mem[3520] = 206;
razn_w_mem[3521] = 206;
razn_w_mem[3522] = 206;
razn_w_mem[3523] = 206;
razn_w_mem[3524] = 206;
razn_w_mem[3525] = 206;
razn_w_mem[3526] = 206;
razn_w_mem[3527] = 206;
razn_w_mem[3528] = 206;
razn_w_mem[3529] = 206;
razn_w_mem[3530] = 206;
razn_w_mem[3531] = 206;
razn_w_mem[3532] = 206;
razn_w_mem[3533] = 206;
razn_w_mem[3534] = 206;
razn_w_mem[3535] = 206;
razn_w_mem[3536] = 206;
razn_w_mem[3537] = 206;
razn_w_mem[3538] = 206;
razn_w_mem[3539] = 206;
razn_w_mem[3540] = 206;
razn_w_mem[3541] = 206;
razn_w_mem[3542] = 206;
razn_w_mem[3543] = 206;
razn_w_mem[3544] = 206;
razn_w_mem[3545] = 206;
razn_w_mem[3546] = 206;
razn_w_mem[3547] = 206;
razn_w_mem[3548] = 206;
razn_w_mem[3549] = 206;
razn_w_mem[3550] = 206;
razn_w_mem[3551] = 206;
razn_w_mem[3552] = 206;
razn_w_mem[3553] = 206;
razn_w_mem[3554] = 206;
razn_w_mem[3555] = 206;
razn_w_mem[3556] = 206;
razn_w_mem[3557] = 206;
razn_w_mem[3558] = 206;
razn_w_mem[3559] = 206;
razn_w_mem[3560] = 206;
razn_w_mem[3561] = 206;
razn_w_mem[3562] = 206;
razn_w_mem[3563] = 206;
razn_w_mem[3564] = 206;
razn_w_mem[3565] = 206;
razn_w_mem[3566] = 206;
razn_w_mem[3567] = 206;
razn_w_mem[3568] = 206;
razn_w_mem[3569] = 206;
razn_w_mem[3570] = 206;
razn_w_mem[3571] = 206;
razn_w_mem[3572] = 206;
razn_w_mem[3573] = 206;
razn_w_mem[3574] = 206;
razn_w_mem[3575] = 206;
razn_w_mem[3576] = 206;
razn_w_mem[3577] = 206;
razn_w_mem[3578] = 206;
razn_w_mem[3579] = 206;
razn_w_mem[3580] = 206;
razn_w_mem[3581] = 206;
razn_w_mem[3582] = 206;
razn_w_mem[3583] = 206;
razn_w_mem[3584] = 176;
razn_w_mem[3585] = 176;
razn_w_mem[3586] = 176;
razn_w_mem[3587] = 176;
razn_w_mem[3588] = 176;
razn_w_mem[3589] = 176;
razn_w_mem[3590] = 176;
razn_w_mem[3591] = 176;
razn_w_mem[3592] = 176;
razn_w_mem[3593] = 176;
razn_w_mem[3594] = 176;
razn_w_mem[3595] = 176;
razn_w_mem[3596] = 176;
razn_w_mem[3597] = 176;
razn_w_mem[3598] = 176;
razn_w_mem[3599] = 176;
razn_w_mem[3600] = 176;
razn_w_mem[3601] = 176;
razn_w_mem[3602] = 176;
razn_w_mem[3603] = 176;
razn_w_mem[3604] = 176;
razn_w_mem[3605] = 176;
razn_w_mem[3606] = 176;
razn_w_mem[3607] = 176;
razn_w_mem[3608] = 176;
razn_w_mem[3609] = 176;
razn_w_mem[3610] = 176;
razn_w_mem[3611] = 176;
razn_w_mem[3612] = 176;
razn_w_mem[3613] = 176;
razn_w_mem[3614] = 176;
razn_w_mem[3615] = 176;
razn_w_mem[3616] = 176;
razn_w_mem[3617] = 176;
razn_w_mem[3618] = 176;
razn_w_mem[3619] = 176;
razn_w_mem[3620] = 176;
razn_w_mem[3621] = 176;
razn_w_mem[3622] = 176;
razn_w_mem[3623] = 176;
razn_w_mem[3624] = 176;
razn_w_mem[3625] = 176;
razn_w_mem[3626] = 176;
razn_w_mem[3627] = 176;
razn_w_mem[3628] = 176;
razn_w_mem[3629] = 176;
razn_w_mem[3630] = 176;
razn_w_mem[3631] = 176;
razn_w_mem[3632] = 176;
razn_w_mem[3633] = 176;
razn_w_mem[3634] = 176;
razn_w_mem[3635] = 176;
razn_w_mem[3636] = 176;
razn_w_mem[3637] = 176;
razn_w_mem[3638] = 176;
razn_w_mem[3639] = 176;
razn_w_mem[3640] = 176;
razn_w_mem[3641] = 176;
razn_w_mem[3642] = 176;
razn_w_mem[3643] = 176;
razn_w_mem[3644] = 176;
razn_w_mem[3645] = 176;
razn_w_mem[3646] = 176;
razn_w_mem[3647] = 176;
razn_w_mem[3648] = 176;
razn_w_mem[3649] = 176;
razn_w_mem[3650] = 176;
razn_w_mem[3651] = 176;
razn_w_mem[3652] = 176;
razn_w_mem[3653] = 176;
razn_w_mem[3654] = 176;
razn_w_mem[3655] = 176;
razn_w_mem[3656] = 176;
razn_w_mem[3657] = 176;
razn_w_mem[3658] = 176;
razn_w_mem[3659] = 176;
razn_w_mem[3660] = 176;
razn_w_mem[3661] = 176;
razn_w_mem[3662] = 176;
razn_w_mem[3663] = 176;
razn_w_mem[3664] = 176;
razn_w_mem[3665] = 176;
razn_w_mem[3666] = 176;
razn_w_mem[3667] = 176;
razn_w_mem[3668] = 176;
razn_w_mem[3669] = 176;
razn_w_mem[3670] = 176;
razn_w_mem[3671] = 176;
razn_w_mem[3672] = 176;
razn_w_mem[3673] = 176;
razn_w_mem[3674] = 176;
razn_w_mem[3675] = 176;
razn_w_mem[3676] = 176;
razn_w_mem[3677] = 176;
razn_w_mem[3678] = 176;
razn_w_mem[3679] = 176;
razn_w_mem[3680] = 176;
razn_w_mem[3681] = 176;
razn_w_mem[3682] = 176;
razn_w_mem[3683] = 176;
razn_w_mem[3684] = 176;
razn_w_mem[3685] = 176;
razn_w_mem[3686] = 176;
razn_w_mem[3687] = 176;
razn_w_mem[3688] = 176;
razn_w_mem[3689] = 176;
razn_w_mem[3690] = 176;
razn_w_mem[3691] = 176;
razn_w_mem[3692] = 176;
razn_w_mem[3693] = 176;
razn_w_mem[3694] = 176;
razn_w_mem[3695] = 176;
razn_w_mem[3696] = 176;
razn_w_mem[3697] = 176;
razn_w_mem[3698] = 176;
razn_w_mem[3699] = 176;
razn_w_mem[3700] = 176;
razn_w_mem[3701] = 176;
razn_w_mem[3702] = 176;
razn_w_mem[3703] = 176;
razn_w_mem[3704] = 176;
razn_w_mem[3705] = 176;
razn_w_mem[3706] = 176;
razn_w_mem[3707] = 176;
razn_w_mem[3708] = 176;
razn_w_mem[3709] = 176;
razn_w_mem[3710] = 176;
razn_w_mem[3711] = 176;
razn_w_mem[3712] = 146;
razn_w_mem[3713] = 146;
razn_w_mem[3714] = 146;
razn_w_mem[3715] = 146;
razn_w_mem[3716] = 146;
razn_w_mem[3717] = 146;
razn_w_mem[3718] = 146;
razn_w_mem[3719] = 146;
razn_w_mem[3720] = 146;
razn_w_mem[3721] = 146;
razn_w_mem[3722] = 146;
razn_w_mem[3723] = 146;
razn_w_mem[3724] = 146;
razn_w_mem[3725] = 146;
razn_w_mem[3726] = 146;
razn_w_mem[3727] = 146;
razn_w_mem[3728] = 146;
razn_w_mem[3729] = 146;
razn_w_mem[3730] = 146;
razn_w_mem[3731] = 146;
razn_w_mem[3732] = 146;
razn_w_mem[3733] = 146;
razn_w_mem[3734] = 146;
razn_w_mem[3735] = 146;
razn_w_mem[3736] = 146;
razn_w_mem[3737] = 146;
razn_w_mem[3738] = 146;
razn_w_mem[3739] = 146;
razn_w_mem[3740] = 146;
razn_w_mem[3741] = 146;
razn_w_mem[3742] = 146;
razn_w_mem[3743] = 146;
razn_w_mem[3744] = 146;
razn_w_mem[3745] = 146;
razn_w_mem[3746] = 146;
razn_w_mem[3747] = 146;
razn_w_mem[3748] = 146;
razn_w_mem[3749] = 146;
razn_w_mem[3750] = 146;
razn_w_mem[3751] = 146;
razn_w_mem[3752] = 146;
razn_w_mem[3753] = 146;
razn_w_mem[3754] = 146;
razn_w_mem[3755] = 146;
razn_w_mem[3756] = 146;
razn_w_mem[3757] = 146;
razn_w_mem[3758] = 146;
razn_w_mem[3759] = 146;
razn_w_mem[3760] = 146;
razn_w_mem[3761] = 146;
razn_w_mem[3762] = 146;
razn_w_mem[3763] = 146;
razn_w_mem[3764] = 146;
razn_w_mem[3765] = 146;
razn_w_mem[3766] = 146;
razn_w_mem[3767] = 146;
razn_w_mem[3768] = 146;
razn_w_mem[3769] = 146;
razn_w_mem[3770] = 146;
razn_w_mem[3771] = 146;
razn_w_mem[3772] = 146;
razn_w_mem[3773] = 146;
razn_w_mem[3774] = 146;
razn_w_mem[3775] = 146;
razn_w_mem[3776] = 146;
razn_w_mem[3777] = 146;
razn_w_mem[3778] = 146;
razn_w_mem[3779] = 146;
razn_w_mem[3780] = 146;
razn_w_mem[3781] = 146;
razn_w_mem[3782] = 146;
razn_w_mem[3783] = 146;
razn_w_mem[3784] = 146;
razn_w_mem[3785] = 146;
razn_w_mem[3786] = 146;
razn_w_mem[3787] = 146;
razn_w_mem[3788] = 146;
razn_w_mem[3789] = 146;
razn_w_mem[3790] = 146;
razn_w_mem[3791] = 146;
razn_w_mem[3792] = 146;
razn_w_mem[3793] = 146;
razn_w_mem[3794] = 146;
razn_w_mem[3795] = 146;
razn_w_mem[3796] = 146;
razn_w_mem[3797] = 146;
razn_w_mem[3798] = 146;
razn_w_mem[3799] = 146;
razn_w_mem[3800] = 146;
razn_w_mem[3801] = 146;
razn_w_mem[3802] = 146;
razn_w_mem[3803] = 146;
razn_w_mem[3804] = 146;
razn_w_mem[3805] = 146;
razn_w_mem[3806] = 146;
razn_w_mem[3807] = 146;
razn_w_mem[3808] = 146;
razn_w_mem[3809] = 146;
razn_w_mem[3810] = 146;
razn_w_mem[3811] = 146;
razn_w_mem[3812] = 146;
razn_w_mem[3813] = 146;
razn_w_mem[3814] = 146;
razn_w_mem[3815] = 146;
razn_w_mem[3816] = 146;
razn_w_mem[3817] = 146;
razn_w_mem[3818] = 146;
razn_w_mem[3819] = 146;
razn_w_mem[3820] = 146;
razn_w_mem[3821] = 146;
razn_w_mem[3822] = 146;
razn_w_mem[3823] = 146;
razn_w_mem[3824] = 146;
razn_w_mem[3825] = 146;
razn_w_mem[3826] = 146;
razn_w_mem[3827] = 146;
razn_w_mem[3828] = 146;
razn_w_mem[3829] = 146;
razn_w_mem[3830] = 146;
razn_w_mem[3831] = 146;
razn_w_mem[3832] = 146;
razn_w_mem[3833] = 146;
razn_w_mem[3834] = 146;
razn_w_mem[3835] = 146;
razn_w_mem[3836] = 146;
razn_w_mem[3837] = 146;
razn_w_mem[3838] = 146;
razn_w_mem[3839] = 146;
razn_w_mem[3840] = 116;
razn_w_mem[3841] = 116;
razn_w_mem[3842] = 116;
razn_w_mem[3843] = 116;
razn_w_mem[3844] = 116;
razn_w_mem[3845] = 116;
razn_w_mem[3846] = 116;
razn_w_mem[3847] = 116;
razn_w_mem[3848] = 116;
razn_w_mem[3849] = 116;
razn_w_mem[3850] = 116;
razn_w_mem[3851] = 116;
razn_w_mem[3852] = 116;
razn_w_mem[3853] = 116;
razn_w_mem[3854] = 116;
razn_w_mem[3855] = 116;
razn_w_mem[3856] = 116;
razn_w_mem[3857] = 116;
razn_w_mem[3858] = 116;
razn_w_mem[3859] = 116;
razn_w_mem[3860] = 116;
razn_w_mem[3861] = 116;
razn_w_mem[3862] = 116;
razn_w_mem[3863] = 116;
razn_w_mem[3864] = 116;
razn_w_mem[3865] = 116;
razn_w_mem[3866] = 116;
razn_w_mem[3867] = 116;
razn_w_mem[3868] = 116;
razn_w_mem[3869] = 116;
razn_w_mem[3870] = 116;
razn_w_mem[3871] = 116;
razn_w_mem[3872] = 116;
razn_w_mem[3873] = 116;
razn_w_mem[3874] = 116;
razn_w_mem[3875] = 116;
razn_w_mem[3876] = 116;
razn_w_mem[3877] = 116;
razn_w_mem[3878] = 116;
razn_w_mem[3879] = 116;
razn_w_mem[3880] = 116;
razn_w_mem[3881] = 116;
razn_w_mem[3882] = 116;
razn_w_mem[3883] = 116;
razn_w_mem[3884] = 116;
razn_w_mem[3885] = 116;
razn_w_mem[3886] = 116;
razn_w_mem[3887] = 116;
razn_w_mem[3888] = 116;
razn_w_mem[3889] = 116;
razn_w_mem[3890] = 116;
razn_w_mem[3891] = 116;
razn_w_mem[3892] = 116;
razn_w_mem[3893] = 116;
razn_w_mem[3894] = 116;
razn_w_mem[3895] = 116;
razn_w_mem[3896] = 116;
razn_w_mem[3897] = 116;
razn_w_mem[3898] = 116;
razn_w_mem[3899] = 116;
razn_w_mem[3900] = 116;
razn_w_mem[3901] = 116;
razn_w_mem[3902] = 116;
razn_w_mem[3903] = 116;
razn_w_mem[3904] = 116;
razn_w_mem[3905] = 116;
razn_w_mem[3906] = 116;
razn_w_mem[3907] = 116;
razn_w_mem[3908] = 116;
razn_w_mem[3909] = 116;
razn_w_mem[3910] = 116;
razn_w_mem[3911] = 116;
razn_w_mem[3912] = 116;
razn_w_mem[3913] = 116;
razn_w_mem[3914] = 116;
razn_w_mem[3915] = 116;
razn_w_mem[3916] = 116;
razn_w_mem[3917] = 116;
razn_w_mem[3918] = 116;
razn_w_mem[3919] = 116;
razn_w_mem[3920] = 116;
razn_w_mem[3921] = 116;
razn_w_mem[3922] = 116;
razn_w_mem[3923] = 116;
razn_w_mem[3924] = 116;
razn_w_mem[3925] = 116;
razn_w_mem[3926] = 116;
razn_w_mem[3927] = 116;
razn_w_mem[3928] = 116;
razn_w_mem[3929] = 116;
razn_w_mem[3930] = 116;
razn_w_mem[3931] = 116;
razn_w_mem[3932] = 116;
razn_w_mem[3933] = 116;
razn_w_mem[3934] = 116;
razn_w_mem[3935] = 116;
razn_w_mem[3936] = 116;
razn_w_mem[3937] = 116;
razn_w_mem[3938] = 116;
razn_w_mem[3939] = 116;
razn_w_mem[3940] = 116;
razn_w_mem[3941] = 116;
razn_w_mem[3942] = 116;
razn_w_mem[3943] = 116;
razn_w_mem[3944] = 116;
razn_w_mem[3945] = 116;
razn_w_mem[3946] = 116;
razn_w_mem[3947] = 116;
razn_w_mem[3948] = 116;
razn_w_mem[3949] = 116;
razn_w_mem[3950] = 116;
razn_w_mem[3951] = 116;
razn_w_mem[3952] = 116;
razn_w_mem[3953] = 116;
razn_w_mem[3954] = 116;
razn_w_mem[3955] = 116;
razn_w_mem[3956] = 116;
razn_w_mem[3957] = 116;
razn_w_mem[3958] = 116;
razn_w_mem[3959] = 116;
razn_w_mem[3960] = 116;
razn_w_mem[3961] = 116;
razn_w_mem[3962] = 116;
razn_w_mem[3963] = 116;
razn_w_mem[3964] = 116;
razn_w_mem[3965] = 116;
razn_w_mem[3966] = 116;
razn_w_mem[3967] = 116;
razn_w_mem[3968] = 86;
razn_w_mem[3969] = 86;
razn_w_mem[3970] = 86;
razn_w_mem[3971] = 86;
razn_w_mem[3972] = 86;
razn_w_mem[3973] = 86;
razn_w_mem[3974] = 86;
razn_w_mem[3975] = 86;
razn_w_mem[3976] = 86;
razn_w_mem[3977] = 86;
razn_w_mem[3978] = 86;
razn_w_mem[3979] = 86;
razn_w_mem[3980] = 86;
razn_w_mem[3981] = 86;
razn_w_mem[3982] = 86;
razn_w_mem[3983] = 86;
razn_w_mem[3984] = 86;
razn_w_mem[3985] = 86;
razn_w_mem[3986] = 86;
razn_w_mem[3987] = 86;
razn_w_mem[3988] = 86;
razn_w_mem[3989] = 86;
razn_w_mem[3990] = 86;
razn_w_mem[3991] = 86;
razn_w_mem[3992] = 86;
razn_w_mem[3993] = 86;
razn_w_mem[3994] = 86;
razn_w_mem[3995] = 86;
razn_w_mem[3996] = 86;
razn_w_mem[3997] = 86;
razn_w_mem[3998] = 86;
razn_w_mem[3999] = 86;
razn_w_mem[4000] = 86;
razn_w_mem[4001] = 86;
razn_w_mem[4002] = 86;
razn_w_mem[4003] = 86;
razn_w_mem[4004] = 86;
razn_w_mem[4005] = 86;
razn_w_mem[4006] = 86;
razn_w_mem[4007] = 86;
razn_w_mem[4008] = 86;
razn_w_mem[4009] = 86;
razn_w_mem[4010] = 86;
razn_w_mem[4011] = 86;
razn_w_mem[4012] = 86;
razn_w_mem[4013] = 86;
razn_w_mem[4014] = 86;
razn_w_mem[4015] = 86;
razn_w_mem[4016] = 86;
razn_w_mem[4017] = 86;
razn_w_mem[4018] = 86;
razn_w_mem[4019] = 86;
razn_w_mem[4020] = 86;
razn_w_mem[4021] = 86;
razn_w_mem[4022] = 86;
razn_w_mem[4023] = 86;
razn_w_mem[4024] = 86;
razn_w_mem[4025] = 86;
razn_w_mem[4026] = 86;
razn_w_mem[4027] = 86;
razn_w_mem[4028] = 86;
razn_w_mem[4029] = 86;
razn_w_mem[4030] = 86;
razn_w_mem[4031] = 86;
razn_w_mem[4032] = 86;
razn_w_mem[4033] = 86;
razn_w_mem[4034] = 86;
razn_w_mem[4035] = 86;
razn_w_mem[4036] = 86;
razn_w_mem[4037] = 86;
razn_w_mem[4038] = 86;
razn_w_mem[4039] = 86;
razn_w_mem[4040] = 86;
razn_w_mem[4041] = 86;
razn_w_mem[4042] = 86;
razn_w_mem[4043] = 86;
razn_w_mem[4044] = 86;
razn_w_mem[4045] = 86;
razn_w_mem[4046] = 86;
razn_w_mem[4047] = 86;
razn_w_mem[4048] = 86;
razn_w_mem[4049] = 86;
razn_w_mem[4050] = 86;
razn_w_mem[4051] = 86;
razn_w_mem[4052] = 86;
razn_w_mem[4053] = 86;
razn_w_mem[4054] = 86;
razn_w_mem[4055] = 86;
razn_w_mem[4056] = 86;
razn_w_mem[4057] = 86;
razn_w_mem[4058] = 86;
razn_w_mem[4059] = 86;
razn_w_mem[4060] = 86;
razn_w_mem[4061] = 86;
razn_w_mem[4062] = 86;
razn_w_mem[4063] = 86;
razn_w_mem[4064] = 86;
razn_w_mem[4065] = 86;
razn_w_mem[4066] = 86;
razn_w_mem[4067] = 86;
razn_w_mem[4068] = 86;
razn_w_mem[4069] = 86;
razn_w_mem[4070] = 86;
razn_w_mem[4071] = 86;
razn_w_mem[4072] = 86;
razn_w_mem[4073] = 86;
razn_w_mem[4074] = 86;
razn_w_mem[4075] = 86;
razn_w_mem[4076] = 86;
razn_w_mem[4077] = 86;
razn_w_mem[4078] = 86;
razn_w_mem[4079] = 86;
razn_w_mem[4080] = 86;
razn_w_mem[4081] = 86;
razn_w_mem[4082] = 86;
razn_w_mem[4083] = 86;
razn_w_mem[4084] = 86;
razn_w_mem[4085] = 86;
razn_w_mem[4086] = 86;
razn_w_mem[4087] = 86;
razn_w_mem[4088] = 86;
razn_w_mem[4089] = 86;
razn_w_mem[4090] = 86;
razn_w_mem[4091] = 86;
razn_w_mem[4092] = 86;
razn_w_mem[4093] = 86;
razn_w_mem[4094] = 86;
razn_w_mem[4095] = 86;
razn_w_mem[4096] = 56;
razn_w_mem[4097] = 56;
razn_w_mem[4098] = 56;
razn_w_mem[4099] = 56;
razn_w_mem[4100] = 56;
razn_w_mem[4101] = 56;
razn_w_mem[4102] = 56;
razn_w_mem[4103] = 56;
razn_w_mem[4104] = 56;
razn_w_mem[4105] = 56;
razn_w_mem[4106] = 56;
razn_w_mem[4107] = 56;
razn_w_mem[4108] = 56;
razn_w_mem[4109] = 56;
razn_w_mem[4110] = 56;
razn_w_mem[4111] = 56;
razn_w_mem[4112] = 56;
razn_w_mem[4113] = 56;
razn_w_mem[4114] = 56;
razn_w_mem[4115] = 56;
razn_w_mem[4116] = 56;
razn_w_mem[4117] = 56;
razn_w_mem[4118] = 56;
razn_w_mem[4119] = 56;
razn_w_mem[4120] = 56;
razn_w_mem[4121] = 56;
razn_w_mem[4122] = 56;
razn_w_mem[4123] = 56;
razn_w_mem[4124] = 56;
razn_w_mem[4125] = 56;
razn_w_mem[4126] = 56;
razn_w_mem[4127] = 56;
razn_w_mem[4128] = 56;
razn_w_mem[4129] = 56;
razn_w_mem[4130] = 56;
razn_w_mem[4131] = 56;
razn_w_mem[4132] = 56;
razn_w_mem[4133] = 56;
razn_w_mem[4134] = 56;
razn_w_mem[4135] = 56;
razn_w_mem[4136] = 56;
razn_w_mem[4137] = 56;
razn_w_mem[4138] = 56;
razn_w_mem[4139] = 56;
razn_w_mem[4140] = 56;
razn_w_mem[4141] = 56;
razn_w_mem[4142] = 56;
razn_w_mem[4143] = 56;
razn_w_mem[4144] = 56;
razn_w_mem[4145] = 56;
razn_w_mem[4146] = 56;
razn_w_mem[4147] = 56;
razn_w_mem[4148] = 56;
razn_w_mem[4149] = 56;
razn_w_mem[4150] = 56;
razn_w_mem[4151] = 56;
razn_w_mem[4152] = 56;
razn_w_mem[4153] = 56;
razn_w_mem[4154] = 56;
razn_w_mem[4155] = 56;
razn_w_mem[4156] = 56;
razn_w_mem[4157] = 56;
razn_w_mem[4158] = 56;
razn_w_mem[4159] = 56;
razn_w_mem[4160] = 56;
razn_w_mem[4161] = 56;
razn_w_mem[4162] = 56;
razn_w_mem[4163] = 56;
razn_w_mem[4164] = 56;
razn_w_mem[4165] = 56;
razn_w_mem[4166] = 56;
razn_w_mem[4167] = 56;
razn_w_mem[4168] = 56;
razn_w_mem[4169] = 56;
razn_w_mem[4170] = 56;
razn_w_mem[4171] = 56;
razn_w_mem[4172] = 56;
razn_w_mem[4173] = 56;
razn_w_mem[4174] = 56;
razn_w_mem[4175] = 56;
razn_w_mem[4176] = 56;
razn_w_mem[4177] = 56;
razn_w_mem[4178] = 56;
razn_w_mem[4179] = 56;
razn_w_mem[4180] = 56;
razn_w_mem[4181] = 56;
razn_w_mem[4182] = 56;
razn_w_mem[4183] = 56;
razn_w_mem[4184] = 56;
razn_w_mem[4185] = 56;
razn_w_mem[4186] = 56;
razn_w_mem[4187] = 56;
razn_w_mem[4188] = 56;
razn_w_mem[4189] = 56;
razn_w_mem[4190] = 56;
razn_w_mem[4191] = 56;
razn_w_mem[4192] = 56;
razn_w_mem[4193] = 56;
razn_w_mem[4194] = 56;
razn_w_mem[4195] = 56;
razn_w_mem[4196] = 56;
razn_w_mem[4197] = 56;
razn_w_mem[4198] = 56;
razn_w_mem[4199] = 56;
razn_w_mem[4200] = 56;
razn_w_mem[4201] = 56;
razn_w_mem[4202] = 56;
razn_w_mem[4203] = 56;
razn_w_mem[4204] = 56;
razn_w_mem[4205] = 56;
razn_w_mem[4206] = 56;
razn_w_mem[4207] = 56;
razn_w_mem[4208] = 56;
razn_w_mem[4209] = 56;
razn_w_mem[4210] = 56;
razn_w_mem[4211] = 56;
razn_w_mem[4212] = 56;
razn_w_mem[4213] = 56;
razn_w_mem[4214] = 56;
razn_w_mem[4215] = 56;
razn_w_mem[4216] = 56;
razn_w_mem[4217] = 56;
razn_w_mem[4218] = 56;
razn_w_mem[4219] = 56;
razn_w_mem[4220] = 56;
razn_w_mem[4221] = 56;
razn_w_mem[4222] = 56;
razn_w_mem[4223] = 56;
razn_w_mem[4224] = 26;
razn_w_mem[4225] = 26;
razn_w_mem[4226] = 26;
razn_w_mem[4227] = 26;
razn_w_mem[4228] = 26;
razn_w_mem[4229] = 26;
razn_w_mem[4230] = 26;
razn_w_mem[4231] = 26;
razn_w_mem[4232] = 26;
razn_w_mem[4233] = 26;
razn_w_mem[4234] = 26;
razn_w_mem[4235] = 26;
razn_w_mem[4236] = 26;
razn_w_mem[4237] = 26;
razn_w_mem[4238] = 26;
razn_w_mem[4239] = 26;
razn_w_mem[4240] = 26;
razn_w_mem[4241] = 26;
razn_w_mem[4242] = 26;
razn_w_mem[4243] = 26;
razn_w_mem[4244] = 26;
razn_w_mem[4245] = 26;
razn_w_mem[4246] = 26;
razn_w_mem[4247] = 26;
razn_w_mem[4248] = 26;
razn_w_mem[4249] = 26;
razn_w_mem[4250] = 26;
razn_w_mem[4251] = 26;
razn_w_mem[4252] = 26;
razn_w_mem[4253] = 26;
razn_w_mem[4254] = 26;
razn_w_mem[4255] = 26;
razn_w_mem[4256] = 26;
razn_w_mem[4257] = 26;
razn_w_mem[4258] = 26;
razn_w_mem[4259] = 26;
razn_w_mem[4260] = 26;
razn_w_mem[4261] = 26;
razn_w_mem[4262] = 26;
razn_w_mem[4263] = 26;
razn_w_mem[4264] = 26;
razn_w_mem[4265] = 26;
razn_w_mem[4266] = 26;
razn_w_mem[4267] = 26;
razn_w_mem[4268] = 26;
razn_w_mem[4269] = 26;
razn_w_mem[4270] = 26;
razn_w_mem[4271] = 26;
razn_w_mem[4272] = 26;
razn_w_mem[4273] = 26;
razn_w_mem[4274] = 26;
razn_w_mem[4275] = 26;
razn_w_mem[4276] = 26;
razn_w_mem[4277] = 26;
razn_w_mem[4278] = 26;
razn_w_mem[4279] = 26;
razn_w_mem[4280] = 26;
razn_w_mem[4281] = 26;
razn_w_mem[4282] = 26;
razn_w_mem[4283] = 26;
razn_w_mem[4284] = 26;
razn_w_mem[4285] = 26;
razn_w_mem[4286] = 26;
razn_w_mem[4287] = 26;
razn_w_mem[4288] = 26;
razn_w_mem[4289] = 26;
razn_w_mem[4290] = 26;
razn_w_mem[4291] = 26;
razn_w_mem[4292] = 26;
razn_w_mem[4293] = 26;
razn_w_mem[4294] = 26;
razn_w_mem[4295] = 26;
razn_w_mem[4296] = 26;
razn_w_mem[4297] = 26;
razn_w_mem[4298] = 26;
razn_w_mem[4299] = 26;
razn_w_mem[4300] = 26;
razn_w_mem[4301] = 26;
razn_w_mem[4302] = 26;
razn_w_mem[4303] = 26;
razn_w_mem[4304] = 26;
razn_w_mem[4305] = 26;
razn_w_mem[4306] = 26;
razn_w_mem[4307] = 26;
razn_w_mem[4308] = 26;
razn_w_mem[4309] = 26;
razn_w_mem[4310] = 26;
razn_w_mem[4311] = 26;
razn_w_mem[4312] = 26;
razn_w_mem[4313] = 26;
razn_w_mem[4314] = 26;
razn_w_mem[4315] = 26;
razn_w_mem[4316] = 26;
razn_w_mem[4317] = 26;
razn_w_mem[4318] = 26;
razn_w_mem[4319] = 26;
razn_w_mem[4320] = 26;
razn_w_mem[4321] = 26;
razn_w_mem[4322] = 26;
razn_w_mem[4323] = 26;
razn_w_mem[4324] = 26;
razn_w_mem[4325] = 26;
razn_w_mem[4326] = 26;
razn_w_mem[4327] = 26;
razn_w_mem[4328] = 26;
razn_w_mem[4329] = 26;
razn_w_mem[4330] = 26;
razn_w_mem[4331] = 26;
razn_w_mem[4332] = 26;
razn_w_mem[4333] = 26;
razn_w_mem[4334] = 26;
razn_w_mem[4335] = 26;
razn_w_mem[4336] = 26;
razn_w_mem[4337] = 26;
razn_w_mem[4338] = 26;
razn_w_mem[4339] = 26;
razn_w_mem[4340] = 26;
razn_w_mem[4341] = 26;
razn_w_mem[4342] = 26;
razn_w_mem[4343] = 26;
razn_w_mem[4344] = 26;
razn_w_mem[4345] = 26;
razn_w_mem[4346] = 26;
razn_w_mem[4347] = 26;
razn_w_mem[4348] = 26;
razn_w_mem[4349] = 26;
razn_w_mem[4350] = 26;
razn_w_mem[4351] = 26;
razn_w_mem[4352] = 250;
razn_w_mem[4353] = 250;
razn_w_mem[4354] = 250;
razn_w_mem[4355] = 250;
razn_w_mem[4356] = 250;
razn_w_mem[4357] = 250;
razn_w_mem[4358] = 250;
razn_w_mem[4359] = 250;
razn_w_mem[4360] = 250;
razn_w_mem[4361] = 250;
razn_w_mem[4362] = 250;
razn_w_mem[4363] = 250;
razn_w_mem[4364] = 250;
razn_w_mem[4365] = 250;
razn_w_mem[4366] = 250;
razn_w_mem[4367] = 250;
razn_w_mem[4368] = 250;
razn_w_mem[4369] = 250;
razn_w_mem[4370] = 250;
razn_w_mem[4371] = 250;
razn_w_mem[4372] = 250;
razn_w_mem[4373] = 250;
razn_w_mem[4374] = 250;
razn_w_mem[4375] = 250;
razn_w_mem[4376] = 250;
razn_w_mem[4377] = 250;
razn_w_mem[4378] = 250;
razn_w_mem[4379] = 250;
razn_w_mem[4380] = 250;
razn_w_mem[4381] = 250;
razn_w_mem[4382] = 250;
razn_w_mem[4383] = 250;
razn_w_mem[4384] = 250;
razn_w_mem[4385] = 250;
razn_w_mem[4386] = 250;
razn_w_mem[4387] = 250;
razn_w_mem[4388] = 250;
razn_w_mem[4389] = 250;
razn_w_mem[4390] = 250;
razn_w_mem[4391] = 250;
razn_w_mem[4392] = 250;
razn_w_mem[4393] = 250;
razn_w_mem[4394] = 250;
razn_w_mem[4395] = 250;
razn_w_mem[4396] = 250;
razn_w_mem[4397] = 250;
razn_w_mem[4398] = 250;
razn_w_mem[4399] = 250;
razn_w_mem[4400] = 250;
razn_w_mem[4401] = 250;
razn_w_mem[4402] = 250;
razn_w_mem[4403] = 250;
razn_w_mem[4404] = 250;
razn_w_mem[4405] = 250;
razn_w_mem[4406] = 250;
razn_w_mem[4407] = 250;
razn_w_mem[4408] = 250;
razn_w_mem[4409] = 250;
razn_w_mem[4410] = 250;
razn_w_mem[4411] = 250;
razn_w_mem[4412] = 250;
razn_w_mem[4413] = 250;
razn_w_mem[4414] = 250;
razn_w_mem[4415] = 250;
razn_w_mem[4416] = 250;
razn_w_mem[4417] = 250;
razn_w_mem[4418] = 250;
razn_w_mem[4419] = 250;
razn_w_mem[4420] = 250;
razn_w_mem[4421] = 250;
razn_w_mem[4422] = 250;
razn_w_mem[4423] = 250;
razn_w_mem[4424] = 250;
razn_w_mem[4425] = 250;
razn_w_mem[4426] = 250;
razn_w_mem[4427] = 250;
razn_w_mem[4428] = 250;
razn_w_mem[4429] = 250;
razn_w_mem[4430] = 250;
razn_w_mem[4431] = 250;
razn_w_mem[4432] = 250;
razn_w_mem[4433] = 250;
razn_w_mem[4434] = 250;
razn_w_mem[4435] = 250;
razn_w_mem[4436] = 250;
razn_w_mem[4437] = 250;
razn_w_mem[4438] = 250;
razn_w_mem[4439] = 250;
razn_w_mem[4440] = 250;
razn_w_mem[4441] = 250;
razn_w_mem[4442] = 250;
razn_w_mem[4443] = 250;
razn_w_mem[4444] = 250;
razn_w_mem[4445] = 250;
razn_w_mem[4446] = 250;
razn_w_mem[4447] = 250;
razn_w_mem[4448] = 250;
razn_w_mem[4449] = 250;
razn_w_mem[4450] = 250;
razn_w_mem[4451] = 250;
razn_w_mem[4452] = 250;
razn_w_mem[4453] = 250;
razn_w_mem[4454] = 250;
razn_w_mem[4455] = 250;
razn_w_mem[4456] = 250;
razn_w_mem[4457] = 250;
razn_w_mem[4458] = 250;
razn_w_mem[4459] = 250;
razn_w_mem[4460] = 250;
razn_w_mem[4461] = 250;
razn_w_mem[4462] = 250;
razn_w_mem[4463] = 250;
razn_w_mem[4464] = 250;
razn_w_mem[4465] = 250;
razn_w_mem[4466] = 250;
razn_w_mem[4467] = 250;
razn_w_mem[4468] = 250;
razn_w_mem[4469] = 250;
razn_w_mem[4470] = 250;
razn_w_mem[4471] = 250;
razn_w_mem[4472] = 250;
razn_w_mem[4473] = 250;
razn_w_mem[4474] = 250;
razn_w_mem[4475] = 250;
razn_w_mem[4476] = 250;
razn_w_mem[4477] = 250;
razn_w_mem[4478] = 250;
razn_w_mem[4479] = 250;
razn_w_mem[4480] = 220;
razn_w_mem[4481] = 220;
razn_w_mem[4482] = 220;
razn_w_mem[4483] = 220;
razn_w_mem[4484] = 220;
razn_w_mem[4485] = 220;
razn_w_mem[4486] = 220;
razn_w_mem[4487] = 220;
razn_w_mem[4488] = 220;
razn_w_mem[4489] = 220;
razn_w_mem[4490] = 220;
razn_w_mem[4491] = 220;
razn_w_mem[4492] = 220;
razn_w_mem[4493] = 220;
razn_w_mem[4494] = 220;
razn_w_mem[4495] = 220;
razn_w_mem[4496] = 220;
razn_w_mem[4497] = 220;
razn_w_mem[4498] = 220;
razn_w_mem[4499] = 220;
razn_w_mem[4500] = 220;
razn_w_mem[4501] = 220;
razn_w_mem[4502] = 220;
razn_w_mem[4503] = 220;
razn_w_mem[4504] = 220;
razn_w_mem[4505] = 220;
razn_w_mem[4506] = 220;
razn_w_mem[4507] = 220;
razn_w_mem[4508] = 220;
razn_w_mem[4509] = 220;
razn_w_mem[4510] = 220;
razn_w_mem[4511] = 220;
razn_w_mem[4512] = 220;
razn_w_mem[4513] = 220;
razn_w_mem[4514] = 220;
razn_w_mem[4515] = 220;
razn_w_mem[4516] = 220;
razn_w_mem[4517] = 220;
razn_w_mem[4518] = 220;
razn_w_mem[4519] = 220;
razn_w_mem[4520] = 220;
razn_w_mem[4521] = 220;
razn_w_mem[4522] = 220;
razn_w_mem[4523] = 220;
razn_w_mem[4524] = 220;
razn_w_mem[4525] = 220;
razn_w_mem[4526] = 220;
razn_w_mem[4527] = 220;
razn_w_mem[4528] = 220;
razn_w_mem[4529] = 220;
razn_w_mem[4530] = 220;
razn_w_mem[4531] = 220;
razn_w_mem[4532] = 220;
razn_w_mem[4533] = 220;
razn_w_mem[4534] = 220;
razn_w_mem[4535] = 220;
razn_w_mem[4536] = 220;
razn_w_mem[4537] = 220;
razn_w_mem[4538] = 220;
razn_w_mem[4539] = 220;
razn_w_mem[4540] = 220;
razn_w_mem[4541] = 220;
razn_w_mem[4542] = 220;
razn_w_mem[4543] = 220;
razn_w_mem[4544] = 220;
razn_w_mem[4545] = 220;
razn_w_mem[4546] = 220;
razn_w_mem[4547] = 220;
razn_w_mem[4548] = 220;
razn_w_mem[4549] = 220;
razn_w_mem[4550] = 220;
razn_w_mem[4551] = 220;
razn_w_mem[4552] = 220;
razn_w_mem[4553] = 220;
razn_w_mem[4554] = 220;
razn_w_mem[4555] = 220;
razn_w_mem[4556] = 220;
razn_w_mem[4557] = 220;
razn_w_mem[4558] = 220;
razn_w_mem[4559] = 220;
razn_w_mem[4560] = 220;
razn_w_mem[4561] = 220;
razn_w_mem[4562] = 220;
razn_w_mem[4563] = 220;
razn_w_mem[4564] = 220;
razn_w_mem[4565] = 220;
razn_w_mem[4566] = 220;
razn_w_mem[4567] = 220;
razn_w_mem[4568] = 220;
razn_w_mem[4569] = 220;
razn_w_mem[4570] = 220;
razn_w_mem[4571] = 220;
razn_w_mem[4572] = 220;
razn_w_mem[4573] = 220;
razn_w_mem[4574] = 220;
razn_w_mem[4575] = 220;
razn_w_mem[4576] = 220;
razn_w_mem[4577] = 220;
razn_w_mem[4578] = 220;
razn_w_mem[4579] = 220;
razn_w_mem[4580] = 220;
razn_w_mem[4581] = 220;
razn_w_mem[4582] = 220;
razn_w_mem[4583] = 220;
razn_w_mem[4584] = 220;
razn_w_mem[4585] = 220;
razn_w_mem[4586] = 220;
razn_w_mem[4587] = 220;
razn_w_mem[4588] = 220;
razn_w_mem[4589] = 220;
razn_w_mem[4590] = 220;
razn_w_mem[4591] = 220;
razn_w_mem[4592] = 220;
razn_w_mem[4593] = 220;
razn_w_mem[4594] = 220;
razn_w_mem[4595] = 220;
razn_w_mem[4596] = 220;
razn_w_mem[4597] = 220;
razn_w_mem[4598] = 220;
razn_w_mem[4599] = 220;
razn_w_mem[4600] = 220;
razn_w_mem[4601] = 220;
razn_w_mem[4602] = 220;
razn_w_mem[4603] = 220;
razn_w_mem[4604] = 220;
razn_w_mem[4605] = 220;
razn_w_mem[4606] = 220;
razn_w_mem[4607] = 220;
razn_w_mem[4608] = 190;
razn_w_mem[4609] = 190;
razn_w_mem[4610] = 190;
razn_w_mem[4611] = 190;
razn_w_mem[4612] = 190;
razn_w_mem[4613] = 190;
razn_w_mem[4614] = 190;
razn_w_mem[4615] = 190;
razn_w_mem[4616] = 190;
razn_w_mem[4617] = 190;
razn_w_mem[4618] = 190;
razn_w_mem[4619] = 190;
razn_w_mem[4620] = 190;
razn_w_mem[4621] = 190;
razn_w_mem[4622] = 190;
razn_w_mem[4623] = 190;
razn_w_mem[4624] = 190;
razn_w_mem[4625] = 190;
razn_w_mem[4626] = 190;
razn_w_mem[4627] = 190;
razn_w_mem[4628] = 190;
razn_w_mem[4629] = 190;
razn_w_mem[4630] = 190;
razn_w_mem[4631] = 190;
razn_w_mem[4632] = 190;
razn_w_mem[4633] = 190;
razn_w_mem[4634] = 190;
razn_w_mem[4635] = 190;
razn_w_mem[4636] = 190;
razn_w_mem[4637] = 190;
razn_w_mem[4638] = 190;
razn_w_mem[4639] = 190;
razn_w_mem[4640] = 190;
razn_w_mem[4641] = 190;
razn_w_mem[4642] = 190;
razn_w_mem[4643] = 190;
razn_w_mem[4644] = 190;
razn_w_mem[4645] = 190;
razn_w_mem[4646] = 190;
razn_w_mem[4647] = 190;
razn_w_mem[4648] = 190;
razn_w_mem[4649] = 190;
razn_w_mem[4650] = 190;
razn_w_mem[4651] = 190;
razn_w_mem[4652] = 190;
razn_w_mem[4653] = 190;
razn_w_mem[4654] = 190;
razn_w_mem[4655] = 190;
razn_w_mem[4656] = 190;
razn_w_mem[4657] = 190;
razn_w_mem[4658] = 190;
razn_w_mem[4659] = 190;
razn_w_mem[4660] = 190;
razn_w_mem[4661] = 190;
razn_w_mem[4662] = 190;
razn_w_mem[4663] = 190;
razn_w_mem[4664] = 190;
razn_w_mem[4665] = 190;
razn_w_mem[4666] = 190;
razn_w_mem[4667] = 190;
razn_w_mem[4668] = 190;
razn_w_mem[4669] = 190;
razn_w_mem[4670] = 190;
razn_w_mem[4671] = 190;
razn_w_mem[4672] = 190;
razn_w_mem[4673] = 190;
razn_w_mem[4674] = 190;
razn_w_mem[4675] = 190;
razn_w_mem[4676] = 190;
razn_w_mem[4677] = 190;
razn_w_mem[4678] = 190;
razn_w_mem[4679] = 190;
razn_w_mem[4680] = 190;
razn_w_mem[4681] = 190;
razn_w_mem[4682] = 190;
razn_w_mem[4683] = 190;
razn_w_mem[4684] = 190;
razn_w_mem[4685] = 190;
razn_w_mem[4686] = 190;
razn_w_mem[4687] = 190;
razn_w_mem[4688] = 190;
razn_w_mem[4689] = 190;
razn_w_mem[4690] = 190;
razn_w_mem[4691] = 190;
razn_w_mem[4692] = 190;
razn_w_mem[4693] = 190;
razn_w_mem[4694] = 190;
razn_w_mem[4695] = 190;
razn_w_mem[4696] = 190;
razn_w_mem[4697] = 190;
razn_w_mem[4698] = 190;
razn_w_mem[4699] = 190;
razn_w_mem[4700] = 190;
razn_w_mem[4701] = 190;
razn_w_mem[4702] = 190;
razn_w_mem[4703] = 190;
razn_w_mem[4704] = 190;
razn_w_mem[4705] = 190;
razn_w_mem[4706] = 190;
razn_w_mem[4707] = 190;
razn_w_mem[4708] = 190;
razn_w_mem[4709] = 190;
razn_w_mem[4710] = 190;
razn_w_mem[4711] = 190;
razn_w_mem[4712] = 190;
razn_w_mem[4713] = 190;
razn_w_mem[4714] = 190;
razn_w_mem[4715] = 190;
razn_w_mem[4716] = 190;
razn_w_mem[4717] = 190;
razn_w_mem[4718] = 190;
razn_w_mem[4719] = 190;
razn_w_mem[4720] = 190;
razn_w_mem[4721] = 190;
razn_w_mem[4722] = 190;
razn_w_mem[4723] = 190;
razn_w_mem[4724] = 190;
razn_w_mem[4725] = 190;
razn_w_mem[4726] = 190;
razn_w_mem[4727] = 190;
razn_w_mem[4728] = 190;
razn_w_mem[4729] = 190;
razn_w_mem[4730] = 190;
razn_w_mem[4731] = 190;
razn_w_mem[4732] = 190;
razn_w_mem[4733] = 190;
razn_w_mem[4734] = 190;
razn_w_mem[4735] = 190;
razn_w_mem[4736] = 160;
razn_w_mem[4737] = 160;
razn_w_mem[4738] = 160;
razn_w_mem[4739] = 160;
razn_w_mem[4740] = 160;
razn_w_mem[4741] = 160;
razn_w_mem[4742] = 160;
razn_w_mem[4743] = 160;
razn_w_mem[4744] = 160;
razn_w_mem[4745] = 160;
razn_w_mem[4746] = 160;
razn_w_mem[4747] = 160;
razn_w_mem[4748] = 160;
razn_w_mem[4749] = 160;
razn_w_mem[4750] = 160;
razn_w_mem[4751] = 160;
razn_w_mem[4752] = 160;
razn_w_mem[4753] = 160;
razn_w_mem[4754] = 160;
razn_w_mem[4755] = 160;
razn_w_mem[4756] = 160;
razn_w_mem[4757] = 160;
razn_w_mem[4758] = 160;
razn_w_mem[4759] = 160;
razn_w_mem[4760] = 160;
razn_w_mem[4761] = 160;
razn_w_mem[4762] = 160;
razn_w_mem[4763] = 160;
razn_w_mem[4764] = 160;
razn_w_mem[4765] = 160;
razn_w_mem[4766] = 160;
razn_w_mem[4767] = 160;
razn_w_mem[4768] = 160;
razn_w_mem[4769] = 160;
razn_w_mem[4770] = 160;
razn_w_mem[4771] = 160;
razn_w_mem[4772] = 160;
razn_w_mem[4773] = 160;
razn_w_mem[4774] = 160;
razn_w_mem[4775] = 160;
razn_w_mem[4776] = 160;
razn_w_mem[4777] = 160;
razn_w_mem[4778] = 160;
razn_w_mem[4779] = 160;
razn_w_mem[4780] = 160;
razn_w_mem[4781] = 160;
razn_w_mem[4782] = 160;
razn_w_mem[4783] = 160;
razn_w_mem[4784] = 160;
razn_w_mem[4785] = 160;
razn_w_mem[4786] = 160;
razn_w_mem[4787] = 160;
razn_w_mem[4788] = 160;
razn_w_mem[4789] = 160;
razn_w_mem[4790] = 160;
razn_w_mem[4791] = 160;
razn_w_mem[4792] = 160;
razn_w_mem[4793] = 160;
razn_w_mem[4794] = 160;
razn_w_mem[4795] = 160;
razn_w_mem[4796] = 160;
razn_w_mem[4797] = 160;
razn_w_mem[4798] = 160;
razn_w_mem[4799] = 160;
razn_w_mem[4800] = 160;
razn_w_mem[4801] = 160;
razn_w_mem[4802] = 160;
razn_w_mem[4803] = 160;
razn_w_mem[4804] = 160;
razn_w_mem[4805] = 160;
razn_w_mem[4806] = 160;
razn_w_mem[4807] = 160;
razn_w_mem[4808] = 160;
razn_w_mem[4809] = 160;
razn_w_mem[4810] = 160;
razn_w_mem[4811] = 160;
razn_w_mem[4812] = 160;
razn_w_mem[4813] = 160;
razn_w_mem[4814] = 160;
razn_w_mem[4815] = 160;
razn_w_mem[4816] = 160;
razn_w_mem[4817] = 160;
razn_w_mem[4818] = 160;
razn_w_mem[4819] = 160;
razn_w_mem[4820] = 160;
razn_w_mem[4821] = 160;
razn_w_mem[4822] = 160;
razn_w_mem[4823] = 160;
razn_w_mem[4824] = 160;
razn_w_mem[4825] = 160;
razn_w_mem[4826] = 160;
razn_w_mem[4827] = 160;
razn_w_mem[4828] = 160;
razn_w_mem[4829] = 160;
razn_w_mem[4830] = 160;
razn_w_mem[4831] = 160;
razn_w_mem[4832] = 160;
razn_w_mem[4833] = 160;
razn_w_mem[4834] = 160;
razn_w_mem[4835] = 160;
razn_w_mem[4836] = 160;
razn_w_mem[4837] = 160;
razn_w_mem[4838] = 160;
razn_w_mem[4839] = 160;
razn_w_mem[4840] = 160;
razn_w_mem[4841] = 160;
razn_w_mem[4842] = 160;
razn_w_mem[4843] = 160;
razn_w_mem[4844] = 160;
razn_w_mem[4845] = 160;
razn_w_mem[4846] = 160;
razn_w_mem[4847] = 160;
razn_w_mem[4848] = 160;
razn_w_mem[4849] = 160;
razn_w_mem[4850] = 160;
razn_w_mem[4851] = 160;
razn_w_mem[4852] = 160;
razn_w_mem[4853] = 160;
razn_w_mem[4854] = 160;
razn_w_mem[4855] = 160;
razn_w_mem[4856] = 160;
razn_w_mem[4857] = 160;
razn_w_mem[4858] = 160;
razn_w_mem[4859] = 160;
razn_w_mem[4860] = 160;
razn_w_mem[4861] = 160;
razn_w_mem[4862] = 160;
razn_w_mem[4863] = 160;
razn_w_mem[4864] = 130;
razn_w_mem[4865] = 130;
razn_w_mem[4866] = 130;
razn_w_mem[4867] = 130;
razn_w_mem[4868] = 130;
razn_w_mem[4869] = 130;
razn_w_mem[4870] = 130;
razn_w_mem[4871] = 130;
razn_w_mem[4872] = 130;
razn_w_mem[4873] = 130;
razn_w_mem[4874] = 130;
razn_w_mem[4875] = 130;
razn_w_mem[4876] = 130;
razn_w_mem[4877] = 130;
razn_w_mem[4878] = 130;
razn_w_mem[4879] = 130;
razn_w_mem[4880] = 130;
razn_w_mem[4881] = 130;
razn_w_mem[4882] = 130;
razn_w_mem[4883] = 130;
razn_w_mem[4884] = 130;
razn_w_mem[4885] = 130;
razn_w_mem[4886] = 130;
razn_w_mem[4887] = 130;
razn_w_mem[4888] = 130;
razn_w_mem[4889] = 130;
razn_w_mem[4890] = 130;
razn_w_mem[4891] = 130;
razn_w_mem[4892] = 130;
razn_w_mem[4893] = 130;
razn_w_mem[4894] = 130;
razn_w_mem[4895] = 130;
razn_w_mem[4896] = 130;
razn_w_mem[4897] = 130;
razn_w_mem[4898] = 130;
razn_w_mem[4899] = 130;
razn_w_mem[4900] = 130;
razn_w_mem[4901] = 130;
razn_w_mem[4902] = 130;
razn_w_mem[4903] = 130;
razn_w_mem[4904] = 130;
razn_w_mem[4905] = 130;
razn_w_mem[4906] = 130;
razn_w_mem[4907] = 130;
razn_w_mem[4908] = 130;
razn_w_mem[4909] = 130;
razn_w_mem[4910] = 130;
razn_w_mem[4911] = 130;
razn_w_mem[4912] = 130;
razn_w_mem[4913] = 130;
razn_w_mem[4914] = 130;
razn_w_mem[4915] = 130;
razn_w_mem[4916] = 130;
razn_w_mem[4917] = 130;
razn_w_mem[4918] = 130;
razn_w_mem[4919] = 130;
razn_w_mem[4920] = 130;
razn_w_mem[4921] = 130;
razn_w_mem[4922] = 130;
razn_w_mem[4923] = 130;
razn_w_mem[4924] = 130;
razn_w_mem[4925] = 130;
razn_w_mem[4926] = 130;
razn_w_mem[4927] = 130;
razn_w_mem[4928] = 130;
razn_w_mem[4929] = 130;
razn_w_mem[4930] = 130;
razn_w_mem[4931] = 130;
razn_w_mem[4932] = 130;
razn_w_mem[4933] = 130;
razn_w_mem[4934] = 130;
razn_w_mem[4935] = 130;
razn_w_mem[4936] = 130;
razn_w_mem[4937] = 130;
razn_w_mem[4938] = 130;
razn_w_mem[4939] = 130;
razn_w_mem[4940] = 130;
razn_w_mem[4941] = 130;
razn_w_mem[4942] = 130;
razn_w_mem[4943] = 130;
razn_w_mem[4944] = 130;
razn_w_mem[4945] = 130;
razn_w_mem[4946] = 130;
razn_w_mem[4947] = 130;
razn_w_mem[4948] = 130;
razn_w_mem[4949] = 130;
razn_w_mem[4950] = 130;
razn_w_mem[4951] = 130;
razn_w_mem[4952] = 130;
razn_w_mem[4953] = 130;
razn_w_mem[4954] = 130;
razn_w_mem[4955] = 130;
razn_w_mem[4956] = 130;
razn_w_mem[4957] = 130;
razn_w_mem[4958] = 130;
razn_w_mem[4959] = 130;
razn_w_mem[4960] = 130;
razn_w_mem[4961] = 130;
razn_w_mem[4962] = 130;
razn_w_mem[4963] = 130;
razn_w_mem[4964] = 130;
razn_w_mem[4965] = 130;
razn_w_mem[4966] = 130;
razn_w_mem[4967] = 130;
razn_w_mem[4968] = 130;
razn_w_mem[4969] = 130;
razn_w_mem[4970] = 130;
razn_w_mem[4971] = 130;
razn_w_mem[4972] = 130;
razn_w_mem[4973] = 130;
razn_w_mem[4974] = 130;
razn_w_mem[4975] = 130;
razn_w_mem[4976] = 130;
razn_w_mem[4977] = 130;
razn_w_mem[4978] = 130;
razn_w_mem[4979] = 130;
razn_w_mem[4980] = 130;
razn_w_mem[4981] = 130;
razn_w_mem[4982] = 130;
razn_w_mem[4983] = 130;
razn_w_mem[4984] = 130;
razn_w_mem[4985] = 130;
razn_w_mem[4986] = 130;
razn_w_mem[4987] = 130;
razn_w_mem[4988] = 130;
razn_w_mem[4989] = 130;
razn_w_mem[4990] = 130;
razn_w_mem[4991] = 130;
razn_w_mem[4992] = 100;
razn_w_mem[4993] = 100;
razn_w_mem[4994] = 100;
razn_w_mem[4995] = 100;
razn_w_mem[4996] = 100;
razn_w_mem[4997] = 100;
razn_w_mem[4998] = 100;
razn_w_mem[4999] = 100;
razn_w_mem[5000] = 100;
razn_w_mem[5001] = 100;
razn_w_mem[5002] = 100;
razn_w_mem[5003] = 100;
razn_w_mem[5004] = 100;
razn_w_mem[5005] = 100;
razn_w_mem[5006] = 100;
razn_w_mem[5007] = 100;
razn_w_mem[5008] = 100;
razn_w_mem[5009] = 100;
razn_w_mem[5010] = 100;
razn_w_mem[5011] = 100;
razn_w_mem[5012] = 100;
razn_w_mem[5013] = 100;
razn_w_mem[5014] = 100;
razn_w_mem[5015] = 100;
razn_w_mem[5016] = 100;
razn_w_mem[5017] = 100;
razn_w_mem[5018] = 100;
razn_w_mem[5019] = 100;
razn_w_mem[5020] = 100;
razn_w_mem[5021] = 100;
razn_w_mem[5022] = 100;
razn_w_mem[5023] = 100;
razn_w_mem[5024] = 100;
razn_w_mem[5025] = 100;
razn_w_mem[5026] = 100;
razn_w_mem[5027] = 100;
razn_w_mem[5028] = 100;
razn_w_mem[5029] = 100;
razn_w_mem[5030] = 100;
razn_w_mem[5031] = 100;
razn_w_mem[5032] = 100;
razn_w_mem[5033] = 100;
razn_w_mem[5034] = 100;
razn_w_mem[5035] = 100;
razn_w_mem[5036] = 100;
razn_w_mem[5037] = 100;
razn_w_mem[5038] = 100;
razn_w_mem[5039] = 100;
razn_w_mem[5040] = 100;
razn_w_mem[5041] = 100;
razn_w_mem[5042] = 100;
razn_w_mem[5043] = 100;
razn_w_mem[5044] = 100;
razn_w_mem[5045] = 100;
razn_w_mem[5046] = 100;
razn_w_mem[5047] = 100;
razn_w_mem[5048] = 100;
razn_w_mem[5049] = 100;
razn_w_mem[5050] = 100;
razn_w_mem[5051] = 100;
razn_w_mem[5052] = 100;
razn_w_mem[5053] = 100;
razn_w_mem[5054] = 100;
razn_w_mem[5055] = 100;
razn_w_mem[5056] = 100;
razn_w_mem[5057] = 100;
razn_w_mem[5058] = 100;
razn_w_mem[5059] = 100;
razn_w_mem[5060] = 100;
razn_w_mem[5061] = 100;
razn_w_mem[5062] = 100;
razn_w_mem[5063] = 100;
razn_w_mem[5064] = 100;
razn_w_mem[5065] = 100;
razn_w_mem[5066] = 100;
razn_w_mem[5067] = 100;
razn_w_mem[5068] = 100;
razn_w_mem[5069] = 100;
razn_w_mem[5070] = 100;
razn_w_mem[5071] = 100;
razn_w_mem[5072] = 100;
razn_w_mem[5073] = 100;
razn_w_mem[5074] = 100;
razn_w_mem[5075] = 100;
razn_w_mem[5076] = 100;
razn_w_mem[5077] = 100;
razn_w_mem[5078] = 100;
razn_w_mem[5079] = 100;
razn_w_mem[5080] = 100;
razn_w_mem[5081] = 100;
razn_w_mem[5082] = 100;
razn_w_mem[5083] = 100;
razn_w_mem[5084] = 100;
razn_w_mem[5085] = 100;
razn_w_mem[5086] = 100;
razn_w_mem[5087] = 100;
razn_w_mem[5088] = 100;
razn_w_mem[5089] = 100;
razn_w_mem[5090] = 100;
razn_w_mem[5091] = 100;
razn_w_mem[5092] = 100;
razn_w_mem[5093] = 100;
razn_w_mem[5094] = 100;
razn_w_mem[5095] = 100;
razn_w_mem[5096] = 100;
razn_w_mem[5097] = 100;
razn_w_mem[5098] = 100;
razn_w_mem[5099] = 100;
razn_w_mem[5100] = 100;
razn_w_mem[5101] = 100;
razn_w_mem[5102] = 100;
razn_w_mem[5103] = 100;
razn_w_mem[5104] = 100;
razn_w_mem[5105] = 100;
razn_w_mem[5106] = 100;
razn_w_mem[5107] = 100;
razn_w_mem[5108] = 100;
razn_w_mem[5109] = 100;
razn_w_mem[5110] = 100;
razn_w_mem[5111] = 100;
razn_w_mem[5112] = 100;
razn_w_mem[5113] = 100;
razn_w_mem[5114] = 100;
razn_w_mem[5115] = 100;
razn_w_mem[5116] = 100;
razn_w_mem[5117] = 100;
razn_w_mem[5118] = 100;
razn_w_mem[5119] = 100;
razn_w_mem[5120] = 70;
razn_w_mem[5121] = 70;
razn_w_mem[5122] = 70;
razn_w_mem[5123] = 70;
razn_w_mem[5124] = 70;
razn_w_mem[5125] = 70;
razn_w_mem[5126] = 70;
razn_w_mem[5127] = 70;
razn_w_mem[5128] = 70;
razn_w_mem[5129] = 70;
razn_w_mem[5130] = 70;
razn_w_mem[5131] = 70;
razn_w_mem[5132] = 70;
razn_w_mem[5133] = 70;
razn_w_mem[5134] = 70;
razn_w_mem[5135] = 70;
razn_w_mem[5136] = 70;
razn_w_mem[5137] = 70;
razn_w_mem[5138] = 70;
razn_w_mem[5139] = 70;
razn_w_mem[5140] = 70;
razn_w_mem[5141] = 70;
razn_w_mem[5142] = 70;
razn_w_mem[5143] = 70;
razn_w_mem[5144] = 70;
razn_w_mem[5145] = 70;
razn_w_mem[5146] = 70;
razn_w_mem[5147] = 70;
razn_w_mem[5148] = 70;
razn_w_mem[5149] = 70;
razn_w_mem[5150] = 70;
razn_w_mem[5151] = 70;
razn_w_mem[5152] = 70;
razn_w_mem[5153] = 70;
razn_w_mem[5154] = 70;
razn_w_mem[5155] = 70;
razn_w_mem[5156] = 70;
razn_w_mem[5157] = 70;
razn_w_mem[5158] = 70;
razn_w_mem[5159] = 70;
razn_w_mem[5160] = 70;
razn_w_mem[5161] = 70;
razn_w_mem[5162] = 70;
razn_w_mem[5163] = 70;
razn_w_mem[5164] = 70;
razn_w_mem[5165] = 70;
razn_w_mem[5166] = 70;
razn_w_mem[5167] = 70;
razn_w_mem[5168] = 70;
razn_w_mem[5169] = 70;
razn_w_mem[5170] = 70;
razn_w_mem[5171] = 70;
razn_w_mem[5172] = 70;
razn_w_mem[5173] = 70;
razn_w_mem[5174] = 70;
razn_w_mem[5175] = 70;
razn_w_mem[5176] = 70;
razn_w_mem[5177] = 70;
razn_w_mem[5178] = 70;
razn_w_mem[5179] = 70;
razn_w_mem[5180] = 70;
razn_w_mem[5181] = 70;
razn_w_mem[5182] = 70;
razn_w_mem[5183] = 70;
razn_w_mem[5184] = 70;
razn_w_mem[5185] = 70;
razn_w_mem[5186] = 70;
razn_w_mem[5187] = 70;
razn_w_mem[5188] = 70;
razn_w_mem[5189] = 70;
razn_w_mem[5190] = 70;
razn_w_mem[5191] = 70;
razn_w_mem[5192] = 70;
razn_w_mem[5193] = 70;
razn_w_mem[5194] = 70;
razn_w_mem[5195] = 70;
razn_w_mem[5196] = 70;
razn_w_mem[5197] = 70;
razn_w_mem[5198] = 70;
razn_w_mem[5199] = 70;
razn_w_mem[5200] = 70;
razn_w_mem[5201] = 70;
razn_w_mem[5202] = 70;
razn_w_mem[5203] = 70;
razn_w_mem[5204] = 70;
razn_w_mem[5205] = 70;
razn_w_mem[5206] = 70;
razn_w_mem[5207] = 70;
razn_w_mem[5208] = 70;
razn_w_mem[5209] = 70;
razn_w_mem[5210] = 70;
razn_w_mem[5211] = 70;
razn_w_mem[5212] = 70;
razn_w_mem[5213] = 70;
razn_w_mem[5214] = 70;
razn_w_mem[5215] = 70;
razn_w_mem[5216] = 70;
razn_w_mem[5217] = 70;
razn_w_mem[5218] = 70;
razn_w_mem[5219] = 70;
razn_w_mem[5220] = 70;
razn_w_mem[5221] = 70;
razn_w_mem[5222] = 70;
razn_w_mem[5223] = 70;
razn_w_mem[5224] = 70;
razn_w_mem[5225] = 70;
razn_w_mem[5226] = 70;
razn_w_mem[5227] = 70;
razn_w_mem[5228] = 70;
razn_w_mem[5229] = 70;
razn_w_mem[5230] = 70;
razn_w_mem[5231] = 70;
razn_w_mem[5232] = 70;
razn_w_mem[5233] = 70;
razn_w_mem[5234] = 70;
razn_w_mem[5235] = 70;
razn_w_mem[5236] = 70;
razn_w_mem[5237] = 70;
razn_w_mem[5238] = 70;
razn_w_mem[5239] = 70;
razn_w_mem[5240] = 70;
razn_w_mem[5241] = 70;
razn_w_mem[5242] = 70;
razn_w_mem[5243] = 70;
razn_w_mem[5244] = 70;
razn_w_mem[5245] = 70;
razn_w_mem[5246] = 70;
razn_w_mem[5247] = 70;
razn_w_mem[5248] = 40;
razn_w_mem[5249] = 40;
razn_w_mem[5250] = 40;
razn_w_mem[5251] = 40;
razn_w_mem[5252] = 40;
razn_w_mem[5253] = 40;
razn_w_mem[5254] = 40;
razn_w_mem[5255] = 40;
razn_w_mem[5256] = 40;
razn_w_mem[5257] = 40;
razn_w_mem[5258] = 40;
razn_w_mem[5259] = 40;
razn_w_mem[5260] = 40;
razn_w_mem[5261] = 40;
razn_w_mem[5262] = 40;
razn_w_mem[5263] = 40;
razn_w_mem[5264] = 40;
razn_w_mem[5265] = 40;
razn_w_mem[5266] = 40;
razn_w_mem[5267] = 40;
razn_w_mem[5268] = 40;
razn_w_mem[5269] = 40;
razn_w_mem[5270] = 40;
razn_w_mem[5271] = 40;
razn_w_mem[5272] = 40;
razn_w_mem[5273] = 40;
razn_w_mem[5274] = 40;
razn_w_mem[5275] = 40;
razn_w_mem[5276] = 40;
razn_w_mem[5277] = 40;
razn_w_mem[5278] = 40;
razn_w_mem[5279] = 40;
razn_w_mem[5280] = 40;
razn_w_mem[5281] = 40;
razn_w_mem[5282] = 40;
razn_w_mem[5283] = 40;
razn_w_mem[5284] = 40;
razn_w_mem[5285] = 40;
razn_w_mem[5286] = 40;
razn_w_mem[5287] = 40;
razn_w_mem[5288] = 40;
razn_w_mem[5289] = 40;
razn_w_mem[5290] = 40;
razn_w_mem[5291] = 40;
razn_w_mem[5292] = 40;
razn_w_mem[5293] = 40;
razn_w_mem[5294] = 40;
razn_w_mem[5295] = 40;
razn_w_mem[5296] = 40;
razn_w_mem[5297] = 40;
razn_w_mem[5298] = 40;
razn_w_mem[5299] = 40;
razn_w_mem[5300] = 40;
razn_w_mem[5301] = 40;
razn_w_mem[5302] = 40;
razn_w_mem[5303] = 40;
razn_w_mem[5304] = 40;
razn_w_mem[5305] = 40;
razn_w_mem[5306] = 40;
razn_w_mem[5307] = 40;
razn_w_mem[5308] = 40;
razn_w_mem[5309] = 40;
razn_w_mem[5310] = 40;
razn_w_mem[5311] = 40;
razn_w_mem[5312] = 40;
razn_w_mem[5313] = 40;
razn_w_mem[5314] = 40;
razn_w_mem[5315] = 40;
razn_w_mem[5316] = 40;
razn_w_mem[5317] = 40;
razn_w_mem[5318] = 40;
razn_w_mem[5319] = 40;
razn_w_mem[5320] = 40;
razn_w_mem[5321] = 40;
razn_w_mem[5322] = 40;
razn_w_mem[5323] = 40;
razn_w_mem[5324] = 40;
razn_w_mem[5325] = 40;
razn_w_mem[5326] = 40;
razn_w_mem[5327] = 40;
razn_w_mem[5328] = 40;
razn_w_mem[5329] = 40;
razn_w_mem[5330] = 40;
razn_w_mem[5331] = 40;
razn_w_mem[5332] = 40;
razn_w_mem[5333] = 40;
razn_w_mem[5334] = 40;
razn_w_mem[5335] = 40;
razn_w_mem[5336] = 40;
razn_w_mem[5337] = 40;
razn_w_mem[5338] = 40;
razn_w_mem[5339] = 40;
razn_w_mem[5340] = 40;
razn_w_mem[5341] = 40;
razn_w_mem[5342] = 40;
razn_w_mem[5343] = 40;
razn_w_mem[5344] = 40;
razn_w_mem[5345] = 40;
razn_w_mem[5346] = 40;
razn_w_mem[5347] = 40;
razn_w_mem[5348] = 40;
razn_w_mem[5349] = 40;
razn_w_mem[5350] = 40;
razn_w_mem[5351] = 40;
razn_w_mem[5352] = 40;
razn_w_mem[5353] = 40;
razn_w_mem[5354] = 40;
razn_w_mem[5355] = 40;
razn_w_mem[5356] = 40;
razn_w_mem[5357] = 40;
razn_w_mem[5358] = 40;
razn_w_mem[5359] = 40;
razn_w_mem[5360] = 40;
razn_w_mem[5361] = 40;
razn_w_mem[5362] = 40;
razn_w_mem[5363] = 40;
razn_w_mem[5364] = 40;
razn_w_mem[5365] = 40;
razn_w_mem[5366] = 40;
razn_w_mem[5367] = 40;
razn_w_mem[5368] = 40;
razn_w_mem[5369] = 40;
razn_w_mem[5370] = 40;
razn_w_mem[5371] = 40;
razn_w_mem[5372] = 40;
razn_w_mem[5373] = 40;
razn_w_mem[5374] = 40;
razn_w_mem[5375] = 40;
razn_w_mem[5376] = 10;
razn_w_mem[5377] = 10;
razn_w_mem[5378] = 10;
razn_w_mem[5379] = 10;
razn_w_mem[5380] = 10;
razn_w_mem[5381] = 10;
razn_w_mem[5382] = 10;
razn_w_mem[5383] = 10;
razn_w_mem[5384] = 10;
razn_w_mem[5385] = 10;
razn_w_mem[5386] = 10;
razn_w_mem[5387] = 10;
razn_w_mem[5388] = 10;
razn_w_mem[5389] = 10;
razn_w_mem[5390] = 10;
razn_w_mem[5391] = 10;
razn_w_mem[5392] = 10;
razn_w_mem[5393] = 10;
razn_w_mem[5394] = 10;
razn_w_mem[5395] = 10;
razn_w_mem[5396] = 10;
razn_w_mem[5397] = 10;
razn_w_mem[5398] = 10;
razn_w_mem[5399] = 10;
razn_w_mem[5400] = 10;
razn_w_mem[5401] = 10;
razn_w_mem[5402] = 10;
razn_w_mem[5403] = 10;
razn_w_mem[5404] = 10;
razn_w_mem[5405] = 10;
razn_w_mem[5406] = 10;
razn_w_mem[5407] = 10;
razn_w_mem[5408] = 10;
razn_w_mem[5409] = 10;
razn_w_mem[5410] = 10;
razn_w_mem[5411] = 10;
razn_w_mem[5412] = 10;
razn_w_mem[5413] = 10;
razn_w_mem[5414] = 10;
razn_w_mem[5415] = 10;
razn_w_mem[5416] = 10;
razn_w_mem[5417] = 10;
razn_w_mem[5418] = 10;
razn_w_mem[5419] = 10;
razn_w_mem[5420] = 10;
razn_w_mem[5421] = 10;
razn_w_mem[5422] = 10;
razn_w_mem[5423] = 10;
razn_w_mem[5424] = 10;
razn_w_mem[5425] = 10;
razn_w_mem[5426] = 10;
razn_w_mem[5427] = 10;
razn_w_mem[5428] = 10;
razn_w_mem[5429] = 10;
razn_w_mem[5430] = 10;
razn_w_mem[5431] = 10;
razn_w_mem[5432] = 10;
razn_w_mem[5433] = 10;
razn_w_mem[5434] = 10;
razn_w_mem[5435] = 10;
razn_w_mem[5436] = 10;
razn_w_mem[5437] = 10;
razn_w_mem[5438] = 10;
razn_w_mem[5439] = 10;
razn_w_mem[5440] = 10;
razn_w_mem[5441] = 10;
razn_w_mem[5442] = 10;
razn_w_mem[5443] = 10;
razn_w_mem[5444] = 10;
razn_w_mem[5445] = 10;
razn_w_mem[5446] = 10;
razn_w_mem[5447] = 10;
razn_w_mem[5448] = 10;
razn_w_mem[5449] = 10;
razn_w_mem[5450] = 10;
razn_w_mem[5451] = 10;
razn_w_mem[5452] = 10;
razn_w_mem[5453] = 10;
razn_w_mem[5454] = 10;
razn_w_mem[5455] = 10;
razn_w_mem[5456] = 10;
razn_w_mem[5457] = 10;
razn_w_mem[5458] = 10;
razn_w_mem[5459] = 10;
razn_w_mem[5460] = 10;
razn_w_mem[5461] = 10;
razn_w_mem[5462] = 10;
razn_w_mem[5463] = 10;
razn_w_mem[5464] = 10;
razn_w_mem[5465] = 10;
razn_w_mem[5466] = 10;
razn_w_mem[5467] = 10;
razn_w_mem[5468] = 10;
razn_w_mem[5469] = 10;
razn_w_mem[5470] = 10;
razn_w_mem[5471] = 10;
razn_w_mem[5472] = 10;
razn_w_mem[5473] = 10;
razn_w_mem[5474] = 10;
razn_w_mem[5475] = 10;
razn_w_mem[5476] = 10;
razn_w_mem[5477] = 10;
razn_w_mem[5478] = 10;
razn_w_mem[5479] = 10;
razn_w_mem[5480] = 10;
razn_w_mem[5481] = 10;
razn_w_mem[5482] = 10;
razn_w_mem[5483] = 10;
razn_w_mem[5484] = 10;
razn_w_mem[5485] = 10;
razn_w_mem[5486] = 10;
razn_w_mem[5487] = 10;
razn_w_mem[5488] = 10;
razn_w_mem[5489] = 10;
razn_w_mem[5490] = 10;
razn_w_mem[5491] = 10;
razn_w_mem[5492] = 10;
razn_w_mem[5493] = 10;
razn_w_mem[5494] = 10;
razn_w_mem[5495] = 10;
razn_w_mem[5496] = 10;
razn_w_mem[5497] = 10;
razn_w_mem[5498] = 10;
razn_w_mem[5499] = 10;
razn_w_mem[5500] = 10;
razn_w_mem[5501] = 10;
razn_w_mem[5502] = 10;
razn_w_mem[5503] = 10;
razn_w_mem[5504] = 234;
razn_w_mem[5505] = 234;
razn_w_mem[5506] = 234;
razn_w_mem[5507] = 234;
razn_w_mem[5508] = 234;
razn_w_mem[5509] = 234;
razn_w_mem[5510] = 234;
razn_w_mem[5511] = 234;
razn_w_mem[5512] = 234;
razn_w_mem[5513] = 234;
razn_w_mem[5514] = 234;
razn_w_mem[5515] = 234;
razn_w_mem[5516] = 234;
razn_w_mem[5517] = 234;
razn_w_mem[5518] = 234;
razn_w_mem[5519] = 234;
razn_w_mem[5520] = 234;
razn_w_mem[5521] = 234;
razn_w_mem[5522] = 234;
razn_w_mem[5523] = 234;
razn_w_mem[5524] = 234;
razn_w_mem[5525] = 234;
razn_w_mem[5526] = 234;
razn_w_mem[5527] = 234;
razn_w_mem[5528] = 234;
razn_w_mem[5529] = 234;
razn_w_mem[5530] = 234;
razn_w_mem[5531] = 234;
razn_w_mem[5532] = 234;
razn_w_mem[5533] = 234;
razn_w_mem[5534] = 234;
razn_w_mem[5535] = 234;
razn_w_mem[5536] = 234;
razn_w_mem[5537] = 234;
razn_w_mem[5538] = 234;
razn_w_mem[5539] = 234;
razn_w_mem[5540] = 234;
razn_w_mem[5541] = 234;
razn_w_mem[5542] = 234;
razn_w_mem[5543] = 234;
razn_w_mem[5544] = 234;
razn_w_mem[5545] = 234;
razn_w_mem[5546] = 234;
razn_w_mem[5547] = 234;
razn_w_mem[5548] = 234;
razn_w_mem[5549] = 234;
razn_w_mem[5550] = 234;
razn_w_mem[5551] = 234;
razn_w_mem[5552] = 234;
razn_w_mem[5553] = 234;
razn_w_mem[5554] = 234;
razn_w_mem[5555] = 234;
razn_w_mem[5556] = 234;
razn_w_mem[5557] = 234;
razn_w_mem[5558] = 234;
razn_w_mem[5559] = 234;
razn_w_mem[5560] = 234;
razn_w_mem[5561] = 234;
razn_w_mem[5562] = 234;
razn_w_mem[5563] = 234;
razn_w_mem[5564] = 234;
razn_w_mem[5565] = 234;
razn_w_mem[5566] = 234;
razn_w_mem[5567] = 234;
razn_w_mem[5568] = 234;
razn_w_mem[5569] = 234;
razn_w_mem[5570] = 234;
razn_w_mem[5571] = 234;
razn_w_mem[5572] = 234;
razn_w_mem[5573] = 234;
razn_w_mem[5574] = 234;
razn_w_mem[5575] = 234;
razn_w_mem[5576] = 234;
razn_w_mem[5577] = 234;
razn_w_mem[5578] = 234;
razn_w_mem[5579] = 234;
razn_w_mem[5580] = 234;
razn_w_mem[5581] = 234;
razn_w_mem[5582] = 234;
razn_w_mem[5583] = 234;
razn_w_mem[5584] = 234;
razn_w_mem[5585] = 234;
razn_w_mem[5586] = 234;
razn_w_mem[5587] = 234;
razn_w_mem[5588] = 234;
razn_w_mem[5589] = 234;
razn_w_mem[5590] = 234;
razn_w_mem[5591] = 234;
razn_w_mem[5592] = 234;
razn_w_mem[5593] = 234;
razn_w_mem[5594] = 234;
razn_w_mem[5595] = 234;
razn_w_mem[5596] = 234;
razn_w_mem[5597] = 234;
razn_w_mem[5598] = 234;
razn_w_mem[5599] = 234;
razn_w_mem[5600] = 234;
razn_w_mem[5601] = 234;
razn_w_mem[5602] = 234;
razn_w_mem[5603] = 234;
razn_w_mem[5604] = 234;
razn_w_mem[5605] = 234;
razn_w_mem[5606] = 234;
razn_w_mem[5607] = 234;
razn_w_mem[5608] = 234;
razn_w_mem[5609] = 234;
razn_w_mem[5610] = 234;
razn_w_mem[5611] = 234;
razn_w_mem[5612] = 234;
razn_w_mem[5613] = 234;
razn_w_mem[5614] = 234;
razn_w_mem[5615] = 234;
razn_w_mem[5616] = 234;
razn_w_mem[5617] = 234;
razn_w_mem[5618] = 234;
razn_w_mem[5619] = 234;
razn_w_mem[5620] = 234;
razn_w_mem[5621] = 234;
razn_w_mem[5622] = 234;
razn_w_mem[5623] = 234;
razn_w_mem[5624] = 234;
razn_w_mem[5625] = 234;
razn_w_mem[5626] = 234;
razn_w_mem[5627] = 234;
razn_w_mem[5628] = 234;
razn_w_mem[5629] = 234;
razn_w_mem[5630] = 234;
razn_w_mem[5631] = 234;
razn_w_mem[5632] = 204;
razn_w_mem[5633] = 204;
razn_w_mem[5634] = 204;
razn_w_mem[5635] = 204;
razn_w_mem[5636] = 204;
razn_w_mem[5637] = 204;
razn_w_mem[5638] = 204;
razn_w_mem[5639] = 204;
razn_w_mem[5640] = 204;
razn_w_mem[5641] = 204;
razn_w_mem[5642] = 204;
razn_w_mem[5643] = 204;
razn_w_mem[5644] = 204;
razn_w_mem[5645] = 204;
razn_w_mem[5646] = 204;
razn_w_mem[5647] = 204;
razn_w_mem[5648] = 204;
razn_w_mem[5649] = 204;
razn_w_mem[5650] = 204;
razn_w_mem[5651] = 204;
razn_w_mem[5652] = 204;
razn_w_mem[5653] = 204;
razn_w_mem[5654] = 204;
razn_w_mem[5655] = 204;
razn_w_mem[5656] = 204;
razn_w_mem[5657] = 204;
razn_w_mem[5658] = 204;
razn_w_mem[5659] = 204;
razn_w_mem[5660] = 204;
razn_w_mem[5661] = 204;
razn_w_mem[5662] = 204;
razn_w_mem[5663] = 204;
razn_w_mem[5664] = 204;
razn_w_mem[5665] = 204;
razn_w_mem[5666] = 204;
razn_w_mem[5667] = 204;
razn_w_mem[5668] = 204;
razn_w_mem[5669] = 204;
razn_w_mem[5670] = 204;
razn_w_mem[5671] = 204;
razn_w_mem[5672] = 204;
razn_w_mem[5673] = 204;
razn_w_mem[5674] = 204;
razn_w_mem[5675] = 204;
razn_w_mem[5676] = 204;
razn_w_mem[5677] = 204;
razn_w_mem[5678] = 204;
razn_w_mem[5679] = 204;
razn_w_mem[5680] = 204;
razn_w_mem[5681] = 204;
razn_w_mem[5682] = 204;
razn_w_mem[5683] = 204;
razn_w_mem[5684] = 204;
razn_w_mem[5685] = 204;
razn_w_mem[5686] = 204;
razn_w_mem[5687] = 204;
razn_w_mem[5688] = 204;
razn_w_mem[5689] = 204;
razn_w_mem[5690] = 204;
razn_w_mem[5691] = 204;
razn_w_mem[5692] = 204;
razn_w_mem[5693] = 204;
razn_w_mem[5694] = 204;
razn_w_mem[5695] = 204;
razn_w_mem[5696] = 204;
razn_w_mem[5697] = 204;
razn_w_mem[5698] = 204;
razn_w_mem[5699] = 204;
razn_w_mem[5700] = 204;
razn_w_mem[5701] = 204;
razn_w_mem[5702] = 204;
razn_w_mem[5703] = 204;
razn_w_mem[5704] = 204;
razn_w_mem[5705] = 204;
razn_w_mem[5706] = 204;
razn_w_mem[5707] = 204;
razn_w_mem[5708] = 204;
razn_w_mem[5709] = 204;
razn_w_mem[5710] = 204;
razn_w_mem[5711] = 204;
razn_w_mem[5712] = 204;
razn_w_mem[5713] = 204;
razn_w_mem[5714] = 204;
razn_w_mem[5715] = 204;
razn_w_mem[5716] = 204;
razn_w_mem[5717] = 204;
razn_w_mem[5718] = 204;
razn_w_mem[5719] = 204;
razn_w_mem[5720] = 204;
razn_w_mem[5721] = 204;
razn_w_mem[5722] = 204;
razn_w_mem[5723] = 204;
razn_w_mem[5724] = 204;
razn_w_mem[5725] = 204;
razn_w_mem[5726] = 204;
razn_w_mem[5727] = 204;
razn_w_mem[5728] = 204;
razn_w_mem[5729] = 204;
razn_w_mem[5730] = 204;
razn_w_mem[5731] = 204;
razn_w_mem[5732] = 204;
razn_w_mem[5733] = 204;
razn_w_mem[5734] = 204;
razn_w_mem[5735] = 204;
razn_w_mem[5736] = 204;
razn_w_mem[5737] = 204;
razn_w_mem[5738] = 204;
razn_w_mem[5739] = 204;
razn_w_mem[5740] = 204;
razn_w_mem[5741] = 204;
razn_w_mem[5742] = 204;
razn_w_mem[5743] = 204;
razn_w_mem[5744] = 204;
razn_w_mem[5745] = 204;
razn_w_mem[5746] = 204;
razn_w_mem[5747] = 204;
razn_w_mem[5748] = 204;
razn_w_mem[5749] = 204;
razn_w_mem[5750] = 204;
razn_w_mem[5751] = 204;
razn_w_mem[5752] = 204;
razn_w_mem[5753] = 204;
razn_w_mem[5754] = 204;
razn_w_mem[5755] = 204;
razn_w_mem[5756] = 204;
razn_w_mem[5757] = 204;
razn_w_mem[5758] = 204;
razn_w_mem[5759] = 204;
razn_w_mem[5760] = 174;
razn_w_mem[5761] = 174;
razn_w_mem[5762] = 174;
razn_w_mem[5763] = 174;
razn_w_mem[5764] = 174;
razn_w_mem[5765] = 174;
razn_w_mem[5766] = 174;
razn_w_mem[5767] = 174;
razn_w_mem[5768] = 174;
razn_w_mem[5769] = 174;
razn_w_mem[5770] = 174;
razn_w_mem[5771] = 174;
razn_w_mem[5772] = 174;
razn_w_mem[5773] = 174;
razn_w_mem[5774] = 174;
razn_w_mem[5775] = 174;
razn_w_mem[5776] = 174;
razn_w_mem[5777] = 174;
razn_w_mem[5778] = 174;
razn_w_mem[5779] = 174;
razn_w_mem[5780] = 174;
razn_w_mem[5781] = 174;
razn_w_mem[5782] = 174;
razn_w_mem[5783] = 174;
razn_w_mem[5784] = 174;
razn_w_mem[5785] = 174;
razn_w_mem[5786] = 174;
razn_w_mem[5787] = 174;
razn_w_mem[5788] = 174;
razn_w_mem[5789] = 174;
razn_w_mem[5790] = 174;
razn_w_mem[5791] = 174;
razn_w_mem[5792] = 174;
razn_w_mem[5793] = 174;
razn_w_mem[5794] = 174;
razn_w_mem[5795] = 174;
razn_w_mem[5796] = 174;
razn_w_mem[5797] = 174;
razn_w_mem[5798] = 174;
razn_w_mem[5799] = 174;
razn_w_mem[5800] = 174;
razn_w_mem[5801] = 174;
razn_w_mem[5802] = 174;
razn_w_mem[5803] = 174;
razn_w_mem[5804] = 174;
razn_w_mem[5805] = 174;
razn_w_mem[5806] = 174;
razn_w_mem[5807] = 174;
razn_w_mem[5808] = 174;
razn_w_mem[5809] = 174;
razn_w_mem[5810] = 174;
razn_w_mem[5811] = 174;
razn_w_mem[5812] = 174;
razn_w_mem[5813] = 174;
razn_w_mem[5814] = 174;
razn_w_mem[5815] = 174;
razn_w_mem[5816] = 174;
razn_w_mem[5817] = 174;
razn_w_mem[5818] = 174;
razn_w_mem[5819] = 174;
razn_w_mem[5820] = 174;
razn_w_mem[5821] = 174;
razn_w_mem[5822] = 174;
razn_w_mem[5823] = 174;
razn_w_mem[5824] = 174;
razn_w_mem[5825] = 174;
razn_w_mem[5826] = 174;
razn_w_mem[5827] = 174;
razn_w_mem[5828] = 174;
razn_w_mem[5829] = 174;
razn_w_mem[5830] = 174;
razn_w_mem[5831] = 174;
razn_w_mem[5832] = 174;
razn_w_mem[5833] = 174;
razn_w_mem[5834] = 174;
razn_w_mem[5835] = 174;
razn_w_mem[5836] = 174;
razn_w_mem[5837] = 174;
razn_w_mem[5838] = 174;
razn_w_mem[5839] = 174;
razn_w_mem[5840] = 174;
razn_w_mem[5841] = 174;
razn_w_mem[5842] = 174;
razn_w_mem[5843] = 174;
razn_w_mem[5844] = 174;
razn_w_mem[5845] = 174;
razn_w_mem[5846] = 174;
razn_w_mem[5847] = 174;
razn_w_mem[5848] = 174;
razn_w_mem[5849] = 174;
razn_w_mem[5850] = 174;
razn_w_mem[5851] = 174;
razn_w_mem[5852] = 174;
razn_w_mem[5853] = 174;
razn_w_mem[5854] = 174;
razn_w_mem[5855] = 174;
razn_w_mem[5856] = 174;
razn_w_mem[5857] = 174;
razn_w_mem[5858] = 174;
razn_w_mem[5859] = 174;
razn_w_mem[5860] = 174;
razn_w_mem[5861] = 174;
razn_w_mem[5862] = 174;
razn_w_mem[5863] = 174;
razn_w_mem[5864] = 174;
razn_w_mem[5865] = 174;
razn_w_mem[5866] = 174;
razn_w_mem[5867] = 174;
razn_w_mem[5868] = 174;
razn_w_mem[5869] = 174;
razn_w_mem[5870] = 174;
razn_w_mem[5871] = 174;
razn_w_mem[5872] = 174;
razn_w_mem[5873] = 174;
razn_w_mem[5874] = 174;
razn_w_mem[5875] = 174;
razn_w_mem[5876] = 174;
razn_w_mem[5877] = 174;
razn_w_mem[5878] = 174;
razn_w_mem[5879] = 174;
razn_w_mem[5880] = 174;
razn_w_mem[5881] = 174;
razn_w_mem[5882] = 174;
razn_w_mem[5883] = 174;
razn_w_mem[5884] = 174;
razn_w_mem[5885] = 174;
razn_w_mem[5886] = 174;
razn_w_mem[5887] = 174;
razn_w_mem[5888] = 144;
razn_w_mem[5889] = 144;
razn_w_mem[5890] = 144;
razn_w_mem[5891] = 144;
razn_w_mem[5892] = 144;
razn_w_mem[5893] = 144;
razn_w_mem[5894] = 144;
razn_w_mem[5895] = 144;
razn_w_mem[5896] = 144;
razn_w_mem[5897] = 144;
razn_w_mem[5898] = 144;
razn_w_mem[5899] = 144;
razn_w_mem[5900] = 144;
razn_w_mem[5901] = 144;
razn_w_mem[5902] = 144;
razn_w_mem[5903] = 144;
razn_w_mem[5904] = 144;
razn_w_mem[5905] = 144;
razn_w_mem[5906] = 144;
razn_w_mem[5907] = 144;
razn_w_mem[5908] = 144;
razn_w_mem[5909] = 144;
razn_w_mem[5910] = 144;
razn_w_mem[5911] = 144;
razn_w_mem[5912] = 144;
razn_w_mem[5913] = 144;
razn_w_mem[5914] = 144;
razn_w_mem[5915] = 144;
razn_w_mem[5916] = 144;
razn_w_mem[5917] = 144;
razn_w_mem[5918] = 144;
razn_w_mem[5919] = 144;
razn_w_mem[5920] = 144;
razn_w_mem[5921] = 144;
razn_w_mem[5922] = 144;
razn_w_mem[5923] = 144;
razn_w_mem[5924] = 144;
razn_w_mem[5925] = 144;
razn_w_mem[5926] = 144;
razn_w_mem[5927] = 144;
razn_w_mem[5928] = 144;
razn_w_mem[5929] = 144;
razn_w_mem[5930] = 144;
razn_w_mem[5931] = 144;
razn_w_mem[5932] = 144;
razn_w_mem[5933] = 144;
razn_w_mem[5934] = 144;
razn_w_mem[5935] = 144;
razn_w_mem[5936] = 144;
razn_w_mem[5937] = 144;
razn_w_mem[5938] = 144;
razn_w_mem[5939] = 144;
razn_w_mem[5940] = 144;
razn_w_mem[5941] = 144;
razn_w_mem[5942] = 144;
razn_w_mem[5943] = 144;
razn_w_mem[5944] = 144;
razn_w_mem[5945] = 144;
razn_w_mem[5946] = 144;
razn_w_mem[5947] = 144;
razn_w_mem[5948] = 144;
razn_w_mem[5949] = 144;
razn_w_mem[5950] = 144;
razn_w_mem[5951] = 144;
razn_w_mem[5952] = 144;
razn_w_mem[5953] = 144;
razn_w_mem[5954] = 144;
razn_w_mem[5955] = 144;
razn_w_mem[5956] = 144;
razn_w_mem[5957] = 144;
razn_w_mem[5958] = 144;
razn_w_mem[5959] = 144;
razn_w_mem[5960] = 144;
razn_w_mem[5961] = 144;
razn_w_mem[5962] = 144;
razn_w_mem[5963] = 144;
razn_w_mem[5964] = 144;
razn_w_mem[5965] = 144;
razn_w_mem[5966] = 144;
razn_w_mem[5967] = 144;
razn_w_mem[5968] = 144;
razn_w_mem[5969] = 144;
razn_w_mem[5970] = 144;
razn_w_mem[5971] = 144;
razn_w_mem[5972] = 144;
razn_w_mem[5973] = 144;
razn_w_mem[5974] = 144;
razn_w_mem[5975] = 144;
razn_w_mem[5976] = 144;
razn_w_mem[5977] = 144;
razn_w_mem[5978] = 144;
razn_w_mem[5979] = 144;
razn_w_mem[5980] = 144;
razn_w_mem[5981] = 144;
razn_w_mem[5982] = 144;
razn_w_mem[5983] = 144;
razn_w_mem[5984] = 144;
razn_w_mem[5985] = 144;
razn_w_mem[5986] = 144;
razn_w_mem[5987] = 144;
razn_w_mem[5988] = 144;
razn_w_mem[5989] = 144;
razn_w_mem[5990] = 144;
razn_w_mem[5991] = 144;
razn_w_mem[5992] = 144;
razn_w_mem[5993] = 144;
razn_w_mem[5994] = 144;
razn_w_mem[5995] = 144;
razn_w_mem[5996] = 144;
razn_w_mem[5997] = 144;
razn_w_mem[5998] = 144;
razn_w_mem[5999] = 144;
razn_w_mem[6000] = 144;
razn_w_mem[6001] = 144;
razn_w_mem[6002] = 144;
razn_w_mem[6003] = 144;
razn_w_mem[6004] = 144;
razn_w_mem[6005] = 144;
razn_w_mem[6006] = 144;
razn_w_mem[6007] = 144;
razn_w_mem[6008] = 144;
razn_w_mem[6009] = 144;
razn_w_mem[6010] = 144;
razn_w_mem[6011] = 144;
razn_w_mem[6012] = 144;
razn_w_mem[6013] = 144;
razn_w_mem[6014] = 144;
razn_w_mem[6015] = 144;
razn_w_mem[6016] = 114;
razn_w_mem[6017] = 114;
razn_w_mem[6018] = 114;
razn_w_mem[6019] = 114;
razn_w_mem[6020] = 114;
razn_w_mem[6021] = 114;
razn_w_mem[6022] = 114;
razn_w_mem[6023] = 114;
razn_w_mem[6024] = 114;
razn_w_mem[6025] = 114;
razn_w_mem[6026] = 114;
razn_w_mem[6027] = 114;
razn_w_mem[6028] = 114;
razn_w_mem[6029] = 114;
razn_w_mem[6030] = 114;
razn_w_mem[6031] = 114;
razn_w_mem[6032] = 114;
razn_w_mem[6033] = 114;
razn_w_mem[6034] = 114;
razn_w_mem[6035] = 114;
razn_w_mem[6036] = 114;
razn_w_mem[6037] = 114;
razn_w_mem[6038] = 114;
razn_w_mem[6039] = 114;
razn_w_mem[6040] = 114;
razn_w_mem[6041] = 114;
razn_w_mem[6042] = 114;
razn_w_mem[6043] = 114;
razn_w_mem[6044] = 114;
razn_w_mem[6045] = 114;
razn_w_mem[6046] = 114;
razn_w_mem[6047] = 114;
razn_w_mem[6048] = 114;
razn_w_mem[6049] = 114;
razn_w_mem[6050] = 114;
razn_w_mem[6051] = 114;
razn_w_mem[6052] = 114;
razn_w_mem[6053] = 114;
razn_w_mem[6054] = 114;
razn_w_mem[6055] = 114;
razn_w_mem[6056] = 114;
razn_w_mem[6057] = 114;
razn_w_mem[6058] = 114;
razn_w_mem[6059] = 114;
razn_w_mem[6060] = 114;
razn_w_mem[6061] = 114;
razn_w_mem[6062] = 114;
razn_w_mem[6063] = 114;
razn_w_mem[6064] = 114;
razn_w_mem[6065] = 114;
razn_w_mem[6066] = 114;
razn_w_mem[6067] = 114;
razn_w_mem[6068] = 114;
razn_w_mem[6069] = 114;
razn_w_mem[6070] = 114;
razn_w_mem[6071] = 114;
razn_w_mem[6072] = 114;
razn_w_mem[6073] = 114;
razn_w_mem[6074] = 114;
razn_w_mem[6075] = 114;
razn_w_mem[6076] = 114;
razn_w_mem[6077] = 114;
razn_w_mem[6078] = 114;
razn_w_mem[6079] = 114;
razn_w_mem[6080] = 114;
razn_w_mem[6081] = 114;
razn_w_mem[6082] = 114;
razn_w_mem[6083] = 114;
razn_w_mem[6084] = 114;
razn_w_mem[6085] = 114;
razn_w_mem[6086] = 114;
razn_w_mem[6087] = 114;
razn_w_mem[6088] = 114;
razn_w_mem[6089] = 114;
razn_w_mem[6090] = 114;
razn_w_mem[6091] = 114;
razn_w_mem[6092] = 114;
razn_w_mem[6093] = 114;
razn_w_mem[6094] = 114;
razn_w_mem[6095] = 114;
razn_w_mem[6096] = 114;
razn_w_mem[6097] = 114;
razn_w_mem[6098] = 114;
razn_w_mem[6099] = 114;
razn_w_mem[6100] = 114;
razn_w_mem[6101] = 114;
razn_w_mem[6102] = 114;
razn_w_mem[6103] = 114;
razn_w_mem[6104] = 114;
razn_w_mem[6105] = 114;
razn_w_mem[6106] = 114;
razn_w_mem[6107] = 114;
razn_w_mem[6108] = 114;
razn_w_mem[6109] = 114;
razn_w_mem[6110] = 114;
razn_w_mem[6111] = 114;
razn_w_mem[6112] = 114;
razn_w_mem[6113] = 114;
razn_w_mem[6114] = 114;
razn_w_mem[6115] = 114;
razn_w_mem[6116] = 114;
razn_w_mem[6117] = 114;
razn_w_mem[6118] = 114;
razn_w_mem[6119] = 114;
razn_w_mem[6120] = 114;
razn_w_mem[6121] = 114;
razn_w_mem[6122] = 114;
razn_w_mem[6123] = 114;
razn_w_mem[6124] = 114;
razn_w_mem[6125] = 114;
razn_w_mem[6126] = 114;
razn_w_mem[6127] = 114;
razn_w_mem[6128] = 114;
razn_w_mem[6129] = 114;
razn_w_mem[6130] = 114;
razn_w_mem[6131] = 114;
razn_w_mem[6132] = 114;
razn_w_mem[6133] = 114;
razn_w_mem[6134] = 114;
razn_w_mem[6135] = 114;
razn_w_mem[6136] = 114;
razn_w_mem[6137] = 114;
razn_w_mem[6138] = 114;
razn_w_mem[6139] = 114;
razn_w_mem[6140] = 114;
razn_w_mem[6141] = 114;
razn_w_mem[6142] = 114;
razn_w_mem[6143] = 114;
razn_w_mem[6144] = 84;
razn_w_mem[6145] = 84;
razn_w_mem[6146] = 84;
razn_w_mem[6147] = 84;
razn_w_mem[6148] = 84;
razn_w_mem[6149] = 84;
razn_w_mem[6150] = 84;
razn_w_mem[6151] = 84;
razn_w_mem[6152] = 84;
razn_w_mem[6153] = 84;
razn_w_mem[6154] = 84;
razn_w_mem[6155] = 84;
razn_w_mem[6156] = 84;
razn_w_mem[6157] = 84;
razn_w_mem[6158] = 84;
razn_w_mem[6159] = 84;
razn_w_mem[6160] = 84;
razn_w_mem[6161] = 84;
razn_w_mem[6162] = 84;
razn_w_mem[6163] = 84;
razn_w_mem[6164] = 84;
razn_w_mem[6165] = 84;
razn_w_mem[6166] = 84;
razn_w_mem[6167] = 84;
razn_w_mem[6168] = 84;
razn_w_mem[6169] = 84;
razn_w_mem[6170] = 84;
razn_w_mem[6171] = 84;
razn_w_mem[6172] = 84;
razn_w_mem[6173] = 84;
razn_w_mem[6174] = 84;
razn_w_mem[6175] = 84;
razn_w_mem[6176] = 84;
razn_w_mem[6177] = 84;
razn_w_mem[6178] = 84;
razn_w_mem[6179] = 84;
razn_w_mem[6180] = 84;
razn_w_mem[6181] = 84;
razn_w_mem[6182] = 84;
razn_w_mem[6183] = 84;
razn_w_mem[6184] = 84;
razn_w_mem[6185] = 84;
razn_w_mem[6186] = 84;
razn_w_mem[6187] = 84;
razn_w_mem[6188] = 84;
razn_w_mem[6189] = 84;
razn_w_mem[6190] = 84;
razn_w_mem[6191] = 84;
razn_w_mem[6192] = 84;
razn_w_mem[6193] = 84;
razn_w_mem[6194] = 84;
razn_w_mem[6195] = 84;
razn_w_mem[6196] = 84;
razn_w_mem[6197] = 84;
razn_w_mem[6198] = 84;
razn_w_mem[6199] = 84;
razn_w_mem[6200] = 84;
razn_w_mem[6201] = 84;
razn_w_mem[6202] = 84;
razn_w_mem[6203] = 84;
razn_w_mem[6204] = 84;
razn_w_mem[6205] = 84;
razn_w_mem[6206] = 84;
razn_w_mem[6207] = 84;
razn_w_mem[6208] = 84;
razn_w_mem[6209] = 84;
razn_w_mem[6210] = 84;
razn_w_mem[6211] = 84;
razn_w_mem[6212] = 84;
razn_w_mem[6213] = 84;
razn_w_mem[6214] = 84;
razn_w_mem[6215] = 84;
razn_w_mem[6216] = 84;
razn_w_mem[6217] = 84;
razn_w_mem[6218] = 84;
razn_w_mem[6219] = 84;
razn_w_mem[6220] = 84;
razn_w_mem[6221] = 84;
razn_w_mem[6222] = 84;
razn_w_mem[6223] = 84;
razn_w_mem[6224] = 84;
razn_w_mem[6225] = 84;
razn_w_mem[6226] = 84;
razn_w_mem[6227] = 84;
razn_w_mem[6228] = 84;
razn_w_mem[6229] = 84;
razn_w_mem[6230] = 84;
razn_w_mem[6231] = 84;
razn_w_mem[6232] = 84;
razn_w_mem[6233] = 84;
razn_w_mem[6234] = 84;
razn_w_mem[6235] = 84;
razn_w_mem[6236] = 84;
razn_w_mem[6237] = 84;
razn_w_mem[6238] = 84;
razn_w_mem[6239] = 84;
razn_w_mem[6240] = 84;
razn_w_mem[6241] = 84;
razn_w_mem[6242] = 84;
razn_w_mem[6243] = 84;
razn_w_mem[6244] = 84;
razn_w_mem[6245] = 84;
razn_w_mem[6246] = 84;
razn_w_mem[6247] = 84;
razn_w_mem[6248] = 84;
razn_w_mem[6249] = 84;
razn_w_mem[6250] = 84;
razn_w_mem[6251] = 84;
razn_w_mem[6252] = 84;
razn_w_mem[6253] = 84;
razn_w_mem[6254] = 84;
razn_w_mem[6255] = 84;
razn_w_mem[6256] = 84;
razn_w_mem[6257] = 84;
razn_w_mem[6258] = 84;
razn_w_mem[6259] = 84;
razn_w_mem[6260] = 84;
razn_w_mem[6261] = 84;
razn_w_mem[6262] = 84;
razn_w_mem[6263] = 84;
razn_w_mem[6264] = 84;
razn_w_mem[6265] = 84;
razn_w_mem[6266] = 84;
razn_w_mem[6267] = 84;
razn_w_mem[6268] = 84;
razn_w_mem[6269] = 84;
razn_w_mem[6270] = 84;
razn_w_mem[6271] = 84;
razn_w_mem[6272] = 54;
razn_w_mem[6273] = 54;
razn_w_mem[6274] = 54;
razn_w_mem[6275] = 54;
razn_w_mem[6276] = 54;
razn_w_mem[6277] = 54;
razn_w_mem[6278] = 54;
razn_w_mem[6279] = 54;
razn_w_mem[6280] = 54;
razn_w_mem[6281] = 54;
razn_w_mem[6282] = 54;
razn_w_mem[6283] = 54;
razn_w_mem[6284] = 54;
razn_w_mem[6285] = 54;
razn_w_mem[6286] = 54;
razn_w_mem[6287] = 54;
razn_w_mem[6288] = 54;
razn_w_mem[6289] = 54;
razn_w_mem[6290] = 54;
razn_w_mem[6291] = 54;
razn_w_mem[6292] = 54;
razn_w_mem[6293] = 54;
razn_w_mem[6294] = 54;
razn_w_mem[6295] = 54;
razn_w_mem[6296] = 54;
razn_w_mem[6297] = 54;
razn_w_mem[6298] = 54;
razn_w_mem[6299] = 54;
razn_w_mem[6300] = 54;
razn_w_mem[6301] = 54;
razn_w_mem[6302] = 54;
razn_w_mem[6303] = 54;
razn_w_mem[6304] = 54;
razn_w_mem[6305] = 54;
razn_w_mem[6306] = 54;
razn_w_mem[6307] = 54;
razn_w_mem[6308] = 54;
razn_w_mem[6309] = 54;
razn_w_mem[6310] = 54;
razn_w_mem[6311] = 54;
razn_w_mem[6312] = 54;
razn_w_mem[6313] = 54;
razn_w_mem[6314] = 54;
razn_w_mem[6315] = 54;
razn_w_mem[6316] = 54;
razn_w_mem[6317] = 54;
razn_w_mem[6318] = 54;
razn_w_mem[6319] = 54;
razn_w_mem[6320] = 54;
razn_w_mem[6321] = 54;
razn_w_mem[6322] = 54;
razn_w_mem[6323] = 54;
razn_w_mem[6324] = 54;
razn_w_mem[6325] = 54;
razn_w_mem[6326] = 54;
razn_w_mem[6327] = 54;
razn_w_mem[6328] = 54;
razn_w_mem[6329] = 54;
razn_w_mem[6330] = 54;
razn_w_mem[6331] = 54;
razn_w_mem[6332] = 54;
razn_w_mem[6333] = 54;
razn_w_mem[6334] = 54;
razn_w_mem[6335] = 54;
razn_w_mem[6336] = 54;
razn_w_mem[6337] = 54;
razn_w_mem[6338] = 54;
razn_w_mem[6339] = 54;
razn_w_mem[6340] = 54;
razn_w_mem[6341] = 54;
razn_w_mem[6342] = 54;
razn_w_mem[6343] = 54;
razn_w_mem[6344] = 54;
razn_w_mem[6345] = 54;
razn_w_mem[6346] = 54;
razn_w_mem[6347] = 54;
razn_w_mem[6348] = 54;
razn_w_mem[6349] = 54;
razn_w_mem[6350] = 54;
razn_w_mem[6351] = 54;
razn_w_mem[6352] = 54;
razn_w_mem[6353] = 54;
razn_w_mem[6354] = 54;
razn_w_mem[6355] = 54;
razn_w_mem[6356] = 54;
razn_w_mem[6357] = 54;
razn_w_mem[6358] = 54;
razn_w_mem[6359] = 54;
razn_w_mem[6360] = 54;
razn_w_mem[6361] = 54;
razn_w_mem[6362] = 54;
razn_w_mem[6363] = 54;
razn_w_mem[6364] = 54;
razn_w_mem[6365] = 54;
razn_w_mem[6366] = 54;
razn_w_mem[6367] = 54;
razn_w_mem[6368] = 54;
razn_w_mem[6369] = 54;
razn_w_mem[6370] = 54;
razn_w_mem[6371] = 54;
razn_w_mem[6372] = 54;
razn_w_mem[6373] = 54;
razn_w_mem[6374] = 54;
razn_w_mem[6375] = 54;
razn_w_mem[6376] = 54;
razn_w_mem[6377] = 54;
razn_w_mem[6378] = 54;
razn_w_mem[6379] = 54;
razn_w_mem[6380] = 54;
razn_w_mem[6381] = 54;
razn_w_mem[6382] = 54;
razn_w_mem[6383] = 54;
razn_w_mem[6384] = 54;
razn_w_mem[6385] = 54;
razn_w_mem[6386] = 54;
razn_w_mem[6387] = 54;
razn_w_mem[6388] = 54;
razn_w_mem[6389] = 54;
razn_w_mem[6390] = 54;
razn_w_mem[6391] = 54;
razn_w_mem[6392] = 54;
razn_w_mem[6393] = 54;
razn_w_mem[6394] = 54;
razn_w_mem[6395] = 54;
razn_w_mem[6396] = 54;
razn_w_mem[6397] = 54;
razn_w_mem[6398] = 54;
razn_w_mem[6399] = 54;
razn_w_mem[6400] = 24;
razn_w_mem[6401] = 24;
razn_w_mem[6402] = 24;
razn_w_mem[6403] = 24;
razn_w_mem[6404] = 24;
razn_w_mem[6405] = 24;
razn_w_mem[6406] = 24;
razn_w_mem[6407] = 24;
razn_w_mem[6408] = 24;
razn_w_mem[6409] = 24;
razn_w_mem[6410] = 24;
razn_w_mem[6411] = 24;
razn_w_mem[6412] = 24;
razn_w_mem[6413] = 24;
razn_w_mem[6414] = 24;
razn_w_mem[6415] = 24;
razn_w_mem[6416] = 24;
razn_w_mem[6417] = 24;
razn_w_mem[6418] = 24;
razn_w_mem[6419] = 24;
razn_w_mem[6420] = 24;
razn_w_mem[6421] = 24;
razn_w_mem[6422] = 24;
razn_w_mem[6423] = 24;
razn_w_mem[6424] = 24;
razn_w_mem[6425] = 24;
razn_w_mem[6426] = 24;
razn_w_mem[6427] = 24;
razn_w_mem[6428] = 24;
razn_w_mem[6429] = 24;
razn_w_mem[6430] = 24;
razn_w_mem[6431] = 24;
razn_w_mem[6432] = 24;
razn_w_mem[6433] = 24;
razn_w_mem[6434] = 24;
razn_w_mem[6435] = 24;
razn_w_mem[6436] = 24;
razn_w_mem[6437] = 24;
razn_w_mem[6438] = 24;
razn_w_mem[6439] = 24;
razn_w_mem[6440] = 24;
razn_w_mem[6441] = 24;
razn_w_mem[6442] = 24;
razn_w_mem[6443] = 24;
razn_w_mem[6444] = 24;
razn_w_mem[6445] = 24;
razn_w_mem[6446] = 24;
razn_w_mem[6447] = 24;
razn_w_mem[6448] = 24;
razn_w_mem[6449] = 24;
razn_w_mem[6450] = 24;
razn_w_mem[6451] = 24;
razn_w_mem[6452] = 24;
razn_w_mem[6453] = 24;
razn_w_mem[6454] = 24;
razn_w_mem[6455] = 24;
razn_w_mem[6456] = 24;
razn_w_mem[6457] = 24;
razn_w_mem[6458] = 24;
razn_w_mem[6459] = 24;
razn_w_mem[6460] = 24;
razn_w_mem[6461] = 24;
razn_w_mem[6462] = 24;
razn_w_mem[6463] = 24;
razn_w_mem[6464] = 24;
razn_w_mem[6465] = 24;
razn_w_mem[6466] = 24;
razn_w_mem[6467] = 24;
razn_w_mem[6468] = 24;
razn_w_mem[6469] = 24;
razn_w_mem[6470] = 24;
razn_w_mem[6471] = 24;
razn_w_mem[6472] = 24;
razn_w_mem[6473] = 24;
razn_w_mem[6474] = 24;
razn_w_mem[6475] = 24;
razn_w_mem[6476] = 24;
razn_w_mem[6477] = 24;
razn_w_mem[6478] = 24;
razn_w_mem[6479] = 24;
razn_w_mem[6480] = 24;
razn_w_mem[6481] = 24;
razn_w_mem[6482] = 24;
razn_w_mem[6483] = 24;
razn_w_mem[6484] = 24;
razn_w_mem[6485] = 24;
razn_w_mem[6486] = 24;
razn_w_mem[6487] = 24;
razn_w_mem[6488] = 24;
razn_w_mem[6489] = 24;
razn_w_mem[6490] = 24;
razn_w_mem[6491] = 24;
razn_w_mem[6492] = 24;
razn_w_mem[6493] = 24;
razn_w_mem[6494] = 24;
razn_w_mem[6495] = 24;
razn_w_mem[6496] = 24;
razn_w_mem[6497] = 24;
razn_w_mem[6498] = 24;
razn_w_mem[6499] = 24;
razn_w_mem[6500] = 24;
razn_w_mem[6501] = 24;
razn_w_mem[6502] = 24;
razn_w_mem[6503] = 24;
razn_w_mem[6504] = 24;
razn_w_mem[6505] = 24;
razn_w_mem[6506] = 24;
razn_w_mem[6507] = 24;
razn_w_mem[6508] = 24;
razn_w_mem[6509] = 24;
razn_w_mem[6510] = 24;
razn_w_mem[6511] = 24;
razn_w_mem[6512] = 24;
razn_w_mem[6513] = 24;
razn_w_mem[6514] = 24;
razn_w_mem[6515] = 24;
razn_w_mem[6516] = 24;
razn_w_mem[6517] = 24;
razn_w_mem[6518] = 24;
razn_w_mem[6519] = 24;
razn_w_mem[6520] = 24;
razn_w_mem[6521] = 24;
razn_w_mem[6522] = 24;
razn_w_mem[6523] = 24;
razn_w_mem[6524] = 24;
razn_w_mem[6525] = 24;
razn_w_mem[6526] = 24;
razn_w_mem[6527] = 24;
razn_w_mem[6528] = 248;
razn_w_mem[6529] = 248;
razn_w_mem[6530] = 248;
razn_w_mem[6531] = 248;
razn_w_mem[6532] = 248;
razn_w_mem[6533] = 248;
razn_w_mem[6534] = 248;
razn_w_mem[6535] = 248;
razn_w_mem[6536] = 248;
razn_w_mem[6537] = 248;
razn_w_mem[6538] = 248;
razn_w_mem[6539] = 248;
razn_w_mem[6540] = 248;
razn_w_mem[6541] = 248;
razn_w_mem[6542] = 248;
razn_w_mem[6543] = 248;
razn_w_mem[6544] = 248;
razn_w_mem[6545] = 248;
razn_w_mem[6546] = 248;
razn_w_mem[6547] = 248;
razn_w_mem[6548] = 248;
razn_w_mem[6549] = 248;
razn_w_mem[6550] = 248;
razn_w_mem[6551] = 248;
razn_w_mem[6552] = 248;
razn_w_mem[6553] = 248;
razn_w_mem[6554] = 248;
razn_w_mem[6555] = 248;
razn_w_mem[6556] = 248;
razn_w_mem[6557] = 248;
razn_w_mem[6558] = 248;
razn_w_mem[6559] = 248;
razn_w_mem[6560] = 248;
razn_w_mem[6561] = 248;
razn_w_mem[6562] = 248;
razn_w_mem[6563] = 248;
razn_w_mem[6564] = 248;
razn_w_mem[6565] = 248;
razn_w_mem[6566] = 248;
razn_w_mem[6567] = 248;
razn_w_mem[6568] = 248;
razn_w_mem[6569] = 248;
razn_w_mem[6570] = 248;
razn_w_mem[6571] = 248;
razn_w_mem[6572] = 248;
razn_w_mem[6573] = 248;
razn_w_mem[6574] = 248;
razn_w_mem[6575] = 248;
razn_w_mem[6576] = 248;
razn_w_mem[6577] = 248;
razn_w_mem[6578] = 248;
razn_w_mem[6579] = 248;
razn_w_mem[6580] = 248;
razn_w_mem[6581] = 248;
razn_w_mem[6582] = 248;
razn_w_mem[6583] = 248;
razn_w_mem[6584] = 248;
razn_w_mem[6585] = 248;
razn_w_mem[6586] = 248;
razn_w_mem[6587] = 248;
razn_w_mem[6588] = 248;
razn_w_mem[6589] = 248;
razn_w_mem[6590] = 248;
razn_w_mem[6591] = 248;
razn_w_mem[6592] = 248;
razn_w_mem[6593] = 248;
razn_w_mem[6594] = 248;
razn_w_mem[6595] = 248;
razn_w_mem[6596] = 248;
razn_w_mem[6597] = 248;
razn_w_mem[6598] = 248;
razn_w_mem[6599] = 248;
razn_w_mem[6600] = 248;
razn_w_mem[6601] = 248;
razn_w_mem[6602] = 248;
razn_w_mem[6603] = 248;
razn_w_mem[6604] = 248;
razn_w_mem[6605] = 248;
razn_w_mem[6606] = 248;
razn_w_mem[6607] = 248;
razn_w_mem[6608] = 248;
razn_w_mem[6609] = 248;
razn_w_mem[6610] = 248;
razn_w_mem[6611] = 248;
razn_w_mem[6612] = 248;
razn_w_mem[6613] = 248;
razn_w_mem[6614] = 248;
razn_w_mem[6615] = 248;
razn_w_mem[6616] = 248;
razn_w_mem[6617] = 248;
razn_w_mem[6618] = 248;
razn_w_mem[6619] = 248;
razn_w_mem[6620] = 248;
razn_w_mem[6621] = 248;
razn_w_mem[6622] = 248;
razn_w_mem[6623] = 248;
razn_w_mem[6624] = 248;
razn_w_mem[6625] = 248;
razn_w_mem[6626] = 248;
razn_w_mem[6627] = 248;
razn_w_mem[6628] = 248;
razn_w_mem[6629] = 248;
razn_w_mem[6630] = 248;
razn_w_mem[6631] = 248;
razn_w_mem[6632] = 248;
razn_w_mem[6633] = 248;
razn_w_mem[6634] = 248;
razn_w_mem[6635] = 248;
razn_w_mem[6636] = 248;
razn_w_mem[6637] = 248;
razn_w_mem[6638] = 248;
razn_w_mem[6639] = 248;
razn_w_mem[6640] = 248;
razn_w_mem[6641] = 248;
razn_w_mem[6642] = 248;
razn_w_mem[6643] = 248;
razn_w_mem[6644] = 248;
razn_w_mem[6645] = 248;
razn_w_mem[6646] = 248;
razn_w_mem[6647] = 248;
razn_w_mem[6648] = 248;
razn_w_mem[6649] = 248;
razn_w_mem[6650] = 248;
razn_w_mem[6651] = 248;
razn_w_mem[6652] = 248;
razn_w_mem[6653] = 248;
razn_w_mem[6654] = 248;
razn_w_mem[6655] = 248;
razn_w_mem[6656] = 218;
razn_w_mem[6657] = 218;
razn_w_mem[6658] = 218;
razn_w_mem[6659] = 218;
razn_w_mem[6660] = 218;
razn_w_mem[6661] = 218;
razn_w_mem[6662] = 218;
razn_w_mem[6663] = 218;
razn_w_mem[6664] = 218;
razn_w_mem[6665] = 218;
razn_w_mem[6666] = 218;
razn_w_mem[6667] = 218;
razn_w_mem[6668] = 218;
razn_w_mem[6669] = 218;
razn_w_mem[6670] = 218;
razn_w_mem[6671] = 218;
razn_w_mem[6672] = 218;
razn_w_mem[6673] = 218;
razn_w_mem[6674] = 218;
razn_w_mem[6675] = 218;
razn_w_mem[6676] = 218;
razn_w_mem[6677] = 218;
razn_w_mem[6678] = 218;
razn_w_mem[6679] = 218;
razn_w_mem[6680] = 218;
razn_w_mem[6681] = 218;
razn_w_mem[6682] = 218;
razn_w_mem[6683] = 218;
razn_w_mem[6684] = 218;
razn_w_mem[6685] = 218;
razn_w_mem[6686] = 218;
razn_w_mem[6687] = 218;
razn_w_mem[6688] = 218;
razn_w_mem[6689] = 218;
razn_w_mem[6690] = 218;
razn_w_mem[6691] = 218;
razn_w_mem[6692] = 218;
razn_w_mem[6693] = 218;
razn_w_mem[6694] = 218;
razn_w_mem[6695] = 218;
razn_w_mem[6696] = 218;
razn_w_mem[6697] = 218;
razn_w_mem[6698] = 218;
razn_w_mem[6699] = 218;
razn_w_mem[6700] = 218;
razn_w_mem[6701] = 218;
razn_w_mem[6702] = 218;
razn_w_mem[6703] = 218;
razn_w_mem[6704] = 218;
razn_w_mem[6705] = 218;
razn_w_mem[6706] = 218;
razn_w_mem[6707] = 218;
razn_w_mem[6708] = 218;
razn_w_mem[6709] = 218;
razn_w_mem[6710] = 218;
razn_w_mem[6711] = 218;
razn_w_mem[6712] = 218;
razn_w_mem[6713] = 218;
razn_w_mem[6714] = 218;
razn_w_mem[6715] = 218;
razn_w_mem[6716] = 218;
razn_w_mem[6717] = 218;
razn_w_mem[6718] = 218;
razn_w_mem[6719] = 218;
razn_w_mem[6720] = 218;
razn_w_mem[6721] = 218;
razn_w_mem[6722] = 218;
razn_w_mem[6723] = 218;
razn_w_mem[6724] = 218;
razn_w_mem[6725] = 218;
razn_w_mem[6726] = 218;
razn_w_mem[6727] = 218;
razn_w_mem[6728] = 218;
razn_w_mem[6729] = 218;
razn_w_mem[6730] = 218;
razn_w_mem[6731] = 218;
razn_w_mem[6732] = 218;
razn_w_mem[6733] = 218;
razn_w_mem[6734] = 218;
razn_w_mem[6735] = 218;
razn_w_mem[6736] = 218;
razn_w_mem[6737] = 218;
razn_w_mem[6738] = 218;
razn_w_mem[6739] = 218;
razn_w_mem[6740] = 218;
razn_w_mem[6741] = 218;
razn_w_mem[6742] = 218;
razn_w_mem[6743] = 218;
razn_w_mem[6744] = 218;
razn_w_mem[6745] = 218;
razn_w_mem[6746] = 218;
razn_w_mem[6747] = 218;
razn_w_mem[6748] = 218;
razn_w_mem[6749] = 218;
razn_w_mem[6750] = 218;
razn_w_mem[6751] = 218;
razn_w_mem[6752] = 218;
razn_w_mem[6753] = 218;
razn_w_mem[6754] = 218;
razn_w_mem[6755] = 218;
razn_w_mem[6756] = 218;
razn_w_mem[6757] = 218;
razn_w_mem[6758] = 218;
razn_w_mem[6759] = 218;
razn_w_mem[6760] = 218;
razn_w_mem[6761] = 218;
razn_w_mem[6762] = 218;
razn_w_mem[6763] = 218;
razn_w_mem[6764] = 218;
razn_w_mem[6765] = 218;
razn_w_mem[6766] = 218;
razn_w_mem[6767] = 218;
razn_w_mem[6768] = 218;
razn_w_mem[6769] = 218;
razn_w_mem[6770] = 218;
razn_w_mem[6771] = 218;
razn_w_mem[6772] = 218;
razn_w_mem[6773] = 218;
razn_w_mem[6774] = 218;
razn_w_mem[6775] = 218;
razn_w_mem[6776] = 218;
razn_w_mem[6777] = 218;
razn_w_mem[6778] = 218;
razn_w_mem[6779] = 218;
razn_w_mem[6780] = 218;
razn_w_mem[6781] = 218;
razn_w_mem[6782] = 218;
razn_w_mem[6783] = 218;
razn_w_mem[6784] = 188;
razn_w_mem[6785] = 188;
razn_w_mem[6786] = 188;
razn_w_mem[6787] = 188;
razn_w_mem[6788] = 188;
razn_w_mem[6789] = 188;
razn_w_mem[6790] = 188;
razn_w_mem[6791] = 188;
razn_w_mem[6792] = 188;
razn_w_mem[6793] = 188;
razn_w_mem[6794] = 188;
razn_w_mem[6795] = 188;
razn_w_mem[6796] = 188;
razn_w_mem[6797] = 188;
razn_w_mem[6798] = 188;
razn_w_mem[6799] = 188;
razn_w_mem[6800] = 188;
razn_w_mem[6801] = 188;
razn_w_mem[6802] = 188;
razn_w_mem[6803] = 188;
razn_w_mem[6804] = 188;
razn_w_mem[6805] = 188;
razn_w_mem[6806] = 188;
razn_w_mem[6807] = 188;
razn_w_mem[6808] = 188;
razn_w_mem[6809] = 188;
razn_w_mem[6810] = 188;
razn_w_mem[6811] = 188;
razn_w_mem[6812] = 188;
razn_w_mem[6813] = 188;
razn_w_mem[6814] = 188;
razn_w_mem[6815] = 188;
razn_w_mem[6816] = 188;
razn_w_mem[6817] = 188;
razn_w_mem[6818] = 188;
razn_w_mem[6819] = 188;
razn_w_mem[6820] = 188;
razn_w_mem[6821] = 188;
razn_w_mem[6822] = 188;
razn_w_mem[6823] = 188;
razn_w_mem[6824] = 188;
razn_w_mem[6825] = 188;
razn_w_mem[6826] = 188;
razn_w_mem[6827] = 188;
razn_w_mem[6828] = 188;
razn_w_mem[6829] = 188;
razn_w_mem[6830] = 188;
razn_w_mem[6831] = 188;
razn_w_mem[6832] = 188;
razn_w_mem[6833] = 188;
razn_w_mem[6834] = 188;
razn_w_mem[6835] = 188;
razn_w_mem[6836] = 188;
razn_w_mem[6837] = 188;
razn_w_mem[6838] = 188;
razn_w_mem[6839] = 188;
razn_w_mem[6840] = 188;
razn_w_mem[6841] = 188;
razn_w_mem[6842] = 188;
razn_w_mem[6843] = 188;
razn_w_mem[6844] = 188;
razn_w_mem[6845] = 188;
razn_w_mem[6846] = 188;
razn_w_mem[6847] = 188;
razn_w_mem[6848] = 188;
razn_w_mem[6849] = 188;
razn_w_mem[6850] = 188;
razn_w_mem[6851] = 188;
razn_w_mem[6852] = 188;
razn_w_mem[6853] = 188;
razn_w_mem[6854] = 188;
razn_w_mem[6855] = 188;
razn_w_mem[6856] = 188;
razn_w_mem[6857] = 188;
razn_w_mem[6858] = 188;
razn_w_mem[6859] = 188;
razn_w_mem[6860] = 188;
razn_w_mem[6861] = 188;
razn_w_mem[6862] = 188;
razn_w_mem[6863] = 188;
razn_w_mem[6864] = 188;
razn_w_mem[6865] = 188;
razn_w_mem[6866] = 188;
razn_w_mem[6867] = 188;
razn_w_mem[6868] = 188;
razn_w_mem[6869] = 188;
razn_w_mem[6870] = 188;
razn_w_mem[6871] = 188;
razn_w_mem[6872] = 188;
razn_w_mem[6873] = 188;
razn_w_mem[6874] = 188;
razn_w_mem[6875] = 188;
razn_w_mem[6876] = 188;
razn_w_mem[6877] = 188;
razn_w_mem[6878] = 188;
razn_w_mem[6879] = 188;
razn_w_mem[6880] = 188;
razn_w_mem[6881] = 188;
razn_w_mem[6882] = 188;
razn_w_mem[6883] = 188;
razn_w_mem[6884] = 188;
razn_w_mem[6885] = 188;
razn_w_mem[6886] = 188;
razn_w_mem[6887] = 188;
razn_w_mem[6888] = 188;
razn_w_mem[6889] = 188;
razn_w_mem[6890] = 188;
razn_w_mem[6891] = 188;
razn_w_mem[6892] = 188;
razn_w_mem[6893] = 188;
razn_w_mem[6894] = 188;
razn_w_mem[6895] = 188;
razn_w_mem[6896] = 188;
razn_w_mem[6897] = 188;
razn_w_mem[6898] = 188;
razn_w_mem[6899] = 188;
razn_w_mem[6900] = 188;
razn_w_mem[6901] = 188;
razn_w_mem[6902] = 188;
razn_w_mem[6903] = 188;
razn_w_mem[6904] = 188;
razn_w_mem[6905] = 188;
razn_w_mem[6906] = 188;
razn_w_mem[6907] = 188;
razn_w_mem[6908] = 188;
razn_w_mem[6909] = 188;
razn_w_mem[6910] = 188;
razn_w_mem[6911] = 188;
razn_w_mem[6912] = 158;
razn_w_mem[6913] = 158;
razn_w_mem[6914] = 158;
razn_w_mem[6915] = 158;
razn_w_mem[6916] = 158;
razn_w_mem[6917] = 158;
razn_w_mem[6918] = 158;
razn_w_mem[6919] = 158;
razn_w_mem[6920] = 158;
razn_w_mem[6921] = 158;
razn_w_mem[6922] = 158;
razn_w_mem[6923] = 158;
razn_w_mem[6924] = 158;
razn_w_mem[6925] = 158;
razn_w_mem[6926] = 158;
razn_w_mem[6927] = 158;
razn_w_mem[6928] = 158;
razn_w_mem[6929] = 158;
razn_w_mem[6930] = 158;
razn_w_mem[6931] = 158;
razn_w_mem[6932] = 158;
razn_w_mem[6933] = 158;
razn_w_mem[6934] = 158;
razn_w_mem[6935] = 158;
razn_w_mem[6936] = 158;
razn_w_mem[6937] = 158;
razn_w_mem[6938] = 158;
razn_w_mem[6939] = 158;
razn_w_mem[6940] = 158;
razn_w_mem[6941] = 158;
razn_w_mem[6942] = 158;
razn_w_mem[6943] = 158;
razn_w_mem[6944] = 158;
razn_w_mem[6945] = 158;
razn_w_mem[6946] = 158;
razn_w_mem[6947] = 158;
razn_w_mem[6948] = 158;
razn_w_mem[6949] = 158;
razn_w_mem[6950] = 158;
razn_w_mem[6951] = 158;
razn_w_mem[6952] = 158;
razn_w_mem[6953] = 158;
razn_w_mem[6954] = 158;
razn_w_mem[6955] = 158;
razn_w_mem[6956] = 158;
razn_w_mem[6957] = 158;
razn_w_mem[6958] = 158;
razn_w_mem[6959] = 158;
razn_w_mem[6960] = 158;
razn_w_mem[6961] = 158;
razn_w_mem[6962] = 158;
razn_w_mem[6963] = 158;
razn_w_mem[6964] = 158;
razn_w_mem[6965] = 158;
razn_w_mem[6966] = 158;
razn_w_mem[6967] = 158;
razn_w_mem[6968] = 158;
razn_w_mem[6969] = 158;
razn_w_mem[6970] = 158;
razn_w_mem[6971] = 158;
razn_w_mem[6972] = 158;
razn_w_mem[6973] = 158;
razn_w_mem[6974] = 158;
razn_w_mem[6975] = 158;
razn_w_mem[6976] = 158;
razn_w_mem[6977] = 158;
razn_w_mem[6978] = 158;
razn_w_mem[6979] = 158;
razn_w_mem[6980] = 158;
razn_w_mem[6981] = 158;
razn_w_mem[6982] = 158;
razn_w_mem[6983] = 158;
razn_w_mem[6984] = 158;
razn_w_mem[6985] = 158;
razn_w_mem[6986] = 158;
razn_w_mem[6987] = 158;
razn_w_mem[6988] = 158;
razn_w_mem[6989] = 158;
razn_w_mem[6990] = 158;
razn_w_mem[6991] = 158;
razn_w_mem[6992] = 158;
razn_w_mem[6993] = 158;
razn_w_mem[6994] = 158;
razn_w_mem[6995] = 158;
razn_w_mem[6996] = 158;
razn_w_mem[6997] = 158;
razn_w_mem[6998] = 158;
razn_w_mem[6999] = 158;
razn_w_mem[7000] = 158;
razn_w_mem[7001] = 158;
razn_w_mem[7002] = 158;
razn_w_mem[7003] = 158;
razn_w_mem[7004] = 158;
razn_w_mem[7005] = 158;
razn_w_mem[7006] = 158;
razn_w_mem[7007] = 158;
razn_w_mem[7008] = 158;
razn_w_mem[7009] = 158;
razn_w_mem[7010] = 158;
razn_w_mem[7011] = 158;
razn_w_mem[7012] = 158;
razn_w_mem[7013] = 158;
razn_w_mem[7014] = 158;
razn_w_mem[7015] = 158;
razn_w_mem[7016] = 158;
razn_w_mem[7017] = 158;
razn_w_mem[7018] = 158;
razn_w_mem[7019] = 158;
razn_w_mem[7020] = 158;
razn_w_mem[7021] = 158;
razn_w_mem[7022] = 158;
razn_w_mem[7023] = 158;
razn_w_mem[7024] = 158;
razn_w_mem[7025] = 158;
razn_w_mem[7026] = 158;
razn_w_mem[7027] = 158;
razn_w_mem[7028] = 158;
razn_w_mem[7029] = 158;
razn_w_mem[7030] = 158;
razn_w_mem[7031] = 158;
razn_w_mem[7032] = 158;
razn_w_mem[7033] = 158;
razn_w_mem[7034] = 158;
razn_w_mem[7035] = 158;
razn_w_mem[7036] = 158;
razn_w_mem[7037] = 158;
razn_w_mem[7038] = 158;
razn_w_mem[7039] = 158;
razn_w_mem[7040] = 128;
razn_w_mem[7041] = 128;
razn_w_mem[7042] = 128;
razn_w_mem[7043] = 128;
razn_w_mem[7044] = 128;
razn_w_mem[7045] = 128;
razn_w_mem[7046] = 128;
razn_w_mem[7047] = 128;
razn_w_mem[7048] = 128;
razn_w_mem[7049] = 128;
razn_w_mem[7050] = 128;
razn_w_mem[7051] = 128;
razn_w_mem[7052] = 128;
razn_w_mem[7053] = 128;
razn_w_mem[7054] = 128;
razn_w_mem[7055] = 128;
razn_w_mem[7056] = 128;
razn_w_mem[7057] = 128;
razn_w_mem[7058] = 128;
razn_w_mem[7059] = 128;
razn_w_mem[7060] = 128;
razn_w_mem[7061] = 128;
razn_w_mem[7062] = 128;
razn_w_mem[7063] = 128;
razn_w_mem[7064] = 128;
razn_w_mem[7065] = 128;
razn_w_mem[7066] = 128;
razn_w_mem[7067] = 128;
razn_w_mem[7068] = 128;
razn_w_mem[7069] = 128;
razn_w_mem[7070] = 128;
razn_w_mem[7071] = 128;
razn_w_mem[7072] = 128;
razn_w_mem[7073] = 128;
razn_w_mem[7074] = 128;
razn_w_mem[7075] = 128;
razn_w_mem[7076] = 128;
razn_w_mem[7077] = 128;
razn_w_mem[7078] = 128;
razn_w_mem[7079] = 128;
razn_w_mem[7080] = 128;
razn_w_mem[7081] = 128;
razn_w_mem[7082] = 128;
razn_w_mem[7083] = 128;
razn_w_mem[7084] = 128;
razn_w_mem[7085] = 128;
razn_w_mem[7086] = 128;
razn_w_mem[7087] = 128;
razn_w_mem[7088] = 128;
razn_w_mem[7089] = 128;
razn_w_mem[7090] = 128;
razn_w_mem[7091] = 128;
razn_w_mem[7092] = 128;
razn_w_mem[7093] = 128;
razn_w_mem[7094] = 128;
razn_w_mem[7095] = 128;
razn_w_mem[7096] = 128;
razn_w_mem[7097] = 128;
razn_w_mem[7098] = 128;
razn_w_mem[7099] = 128;
razn_w_mem[7100] = 128;
razn_w_mem[7101] = 128;
razn_w_mem[7102] = 128;
razn_w_mem[7103] = 128;
razn_w_mem[7104] = 128;
razn_w_mem[7105] = 128;
razn_w_mem[7106] = 128;
razn_w_mem[7107] = 128;
razn_w_mem[7108] = 128;
razn_w_mem[7109] = 128;
razn_w_mem[7110] = 128;
razn_w_mem[7111] = 128;
razn_w_mem[7112] = 128;
razn_w_mem[7113] = 128;
razn_w_mem[7114] = 128;
razn_w_mem[7115] = 128;
razn_w_mem[7116] = 128;
razn_w_mem[7117] = 128;
razn_w_mem[7118] = 128;
razn_w_mem[7119] = 128;
razn_w_mem[7120] = 128;
razn_w_mem[7121] = 128;
razn_w_mem[7122] = 128;
razn_w_mem[7123] = 128;
razn_w_mem[7124] = 128;
razn_w_mem[7125] = 128;
razn_w_mem[7126] = 128;
razn_w_mem[7127] = 128;
razn_w_mem[7128] = 128;
razn_w_mem[7129] = 128;
razn_w_mem[7130] = 128;
razn_w_mem[7131] = 128;
razn_w_mem[7132] = 128;
razn_w_mem[7133] = 128;
razn_w_mem[7134] = 128;
razn_w_mem[7135] = 128;
razn_w_mem[7136] = 128;
razn_w_mem[7137] = 128;
razn_w_mem[7138] = 128;
razn_w_mem[7139] = 128;
razn_w_mem[7140] = 128;
razn_w_mem[7141] = 128;
razn_w_mem[7142] = 128;
razn_w_mem[7143] = 128;
razn_w_mem[7144] = 128;
razn_w_mem[7145] = 128;
razn_w_mem[7146] = 128;
razn_w_mem[7147] = 128;
razn_w_mem[7148] = 128;
razn_w_mem[7149] = 128;
razn_w_mem[7150] = 128;
razn_w_mem[7151] = 128;
razn_w_mem[7152] = 128;
razn_w_mem[7153] = 128;
razn_w_mem[7154] = 128;
razn_w_mem[7155] = 128;
razn_w_mem[7156] = 128;
razn_w_mem[7157] = 128;
razn_w_mem[7158] = 128;
razn_w_mem[7159] = 128;
razn_w_mem[7160] = 128;
razn_w_mem[7161] = 128;
razn_w_mem[7162] = 128;
razn_w_mem[7163] = 128;
razn_w_mem[7164] = 128;
razn_w_mem[7165] = 128;
razn_w_mem[7166] = 128;
razn_w_mem[7167] = 128;
razn_w_mem[7168] = 98;
razn_w_mem[7169] = 98;
razn_w_mem[7170] = 98;
razn_w_mem[7171] = 98;
razn_w_mem[7172] = 98;
razn_w_mem[7173] = 98;
razn_w_mem[7174] = 98;
razn_w_mem[7175] = 98;
razn_w_mem[7176] = 98;
razn_w_mem[7177] = 98;
razn_w_mem[7178] = 98;
razn_w_mem[7179] = 98;
razn_w_mem[7180] = 98;
razn_w_mem[7181] = 98;
razn_w_mem[7182] = 98;
razn_w_mem[7183] = 98;
razn_w_mem[7184] = 98;
razn_w_mem[7185] = 98;
razn_w_mem[7186] = 98;
razn_w_mem[7187] = 98;
razn_w_mem[7188] = 98;
razn_w_mem[7189] = 98;
razn_w_mem[7190] = 98;
razn_w_mem[7191] = 98;
razn_w_mem[7192] = 98;
razn_w_mem[7193] = 98;
razn_w_mem[7194] = 98;
razn_w_mem[7195] = 98;
razn_w_mem[7196] = 98;
razn_w_mem[7197] = 98;
razn_w_mem[7198] = 98;
razn_w_mem[7199] = 98;
razn_w_mem[7200] = 98;
razn_w_mem[7201] = 98;
razn_w_mem[7202] = 98;
razn_w_mem[7203] = 98;
razn_w_mem[7204] = 98;
razn_w_mem[7205] = 98;
razn_w_mem[7206] = 98;
razn_w_mem[7207] = 98;
razn_w_mem[7208] = 98;
razn_w_mem[7209] = 98;
razn_w_mem[7210] = 98;
razn_w_mem[7211] = 98;
razn_w_mem[7212] = 98;
razn_w_mem[7213] = 98;
razn_w_mem[7214] = 98;
razn_w_mem[7215] = 98;
razn_w_mem[7216] = 98;
razn_w_mem[7217] = 98;
razn_w_mem[7218] = 98;
razn_w_mem[7219] = 98;
razn_w_mem[7220] = 98;
razn_w_mem[7221] = 98;
razn_w_mem[7222] = 98;
razn_w_mem[7223] = 98;
razn_w_mem[7224] = 98;
razn_w_mem[7225] = 98;
razn_w_mem[7226] = 98;
razn_w_mem[7227] = 98;
razn_w_mem[7228] = 98;
razn_w_mem[7229] = 98;
razn_w_mem[7230] = 98;
razn_w_mem[7231] = 98;
razn_w_mem[7232] = 98;
razn_w_mem[7233] = 98;
razn_w_mem[7234] = 98;
razn_w_mem[7235] = 98;
razn_w_mem[7236] = 98;
razn_w_mem[7237] = 98;
razn_w_mem[7238] = 98;
razn_w_mem[7239] = 98;
razn_w_mem[7240] = 98;
razn_w_mem[7241] = 98;
razn_w_mem[7242] = 98;
razn_w_mem[7243] = 98;
razn_w_mem[7244] = 98;
razn_w_mem[7245] = 98;
razn_w_mem[7246] = 98;
razn_w_mem[7247] = 98;
razn_w_mem[7248] = 98;
razn_w_mem[7249] = 98;
razn_w_mem[7250] = 98;
razn_w_mem[7251] = 98;
razn_w_mem[7252] = 98;
razn_w_mem[7253] = 98;
razn_w_mem[7254] = 98;
razn_w_mem[7255] = 98;
razn_w_mem[7256] = 98;
razn_w_mem[7257] = 98;
razn_w_mem[7258] = 98;
razn_w_mem[7259] = 98;
razn_w_mem[7260] = 98;
razn_w_mem[7261] = 98;
razn_w_mem[7262] = 98;
razn_w_mem[7263] = 98;
razn_w_mem[7264] = 98;
razn_w_mem[7265] = 98;
razn_w_mem[7266] = 98;
razn_w_mem[7267] = 98;
razn_w_mem[7268] = 98;
razn_w_mem[7269] = 98;
razn_w_mem[7270] = 98;
razn_w_mem[7271] = 98;
razn_w_mem[7272] = 98;
razn_w_mem[7273] = 98;
razn_w_mem[7274] = 98;
razn_w_mem[7275] = 98;
razn_w_mem[7276] = 98;
razn_w_mem[7277] = 98;
razn_w_mem[7278] = 98;
razn_w_mem[7279] = 98;
razn_w_mem[7280] = 98;
razn_w_mem[7281] = 98;
razn_w_mem[7282] = 98;
razn_w_mem[7283] = 98;
razn_w_mem[7284] = 98;
razn_w_mem[7285] = 98;
razn_w_mem[7286] = 98;
razn_w_mem[7287] = 98;
razn_w_mem[7288] = 98;
razn_w_mem[7289] = 98;
razn_w_mem[7290] = 98;
razn_w_mem[7291] = 98;
razn_w_mem[7292] = 98;
razn_w_mem[7293] = 98;
razn_w_mem[7294] = 98;
razn_w_mem[7295] = 98;
razn_w_mem[7296] = 68;
razn_w_mem[7297] = 68;
razn_w_mem[7298] = 68;
razn_w_mem[7299] = 68;
razn_w_mem[7300] = 68;
razn_w_mem[7301] = 68;
razn_w_mem[7302] = 68;
razn_w_mem[7303] = 68;
razn_w_mem[7304] = 68;
razn_w_mem[7305] = 68;
razn_w_mem[7306] = 68;
razn_w_mem[7307] = 68;
razn_w_mem[7308] = 68;
razn_w_mem[7309] = 68;
razn_w_mem[7310] = 68;
razn_w_mem[7311] = 68;
razn_w_mem[7312] = 68;
razn_w_mem[7313] = 68;
razn_w_mem[7314] = 68;
razn_w_mem[7315] = 68;
razn_w_mem[7316] = 68;
razn_w_mem[7317] = 68;
razn_w_mem[7318] = 68;
razn_w_mem[7319] = 68;
razn_w_mem[7320] = 68;
razn_w_mem[7321] = 68;
razn_w_mem[7322] = 68;
razn_w_mem[7323] = 68;
razn_w_mem[7324] = 68;
razn_w_mem[7325] = 68;
razn_w_mem[7326] = 68;
razn_w_mem[7327] = 68;
razn_w_mem[7328] = 68;
razn_w_mem[7329] = 68;
razn_w_mem[7330] = 68;
razn_w_mem[7331] = 68;
razn_w_mem[7332] = 68;
razn_w_mem[7333] = 68;
razn_w_mem[7334] = 68;
razn_w_mem[7335] = 68;
razn_w_mem[7336] = 68;
razn_w_mem[7337] = 68;
razn_w_mem[7338] = 68;
razn_w_mem[7339] = 68;
razn_w_mem[7340] = 68;
razn_w_mem[7341] = 68;
razn_w_mem[7342] = 68;
razn_w_mem[7343] = 68;
razn_w_mem[7344] = 68;
razn_w_mem[7345] = 68;
razn_w_mem[7346] = 68;
razn_w_mem[7347] = 68;
razn_w_mem[7348] = 68;
razn_w_mem[7349] = 68;
razn_w_mem[7350] = 68;
razn_w_mem[7351] = 68;
razn_w_mem[7352] = 68;
razn_w_mem[7353] = 68;
razn_w_mem[7354] = 68;
razn_w_mem[7355] = 68;
razn_w_mem[7356] = 68;
razn_w_mem[7357] = 68;
razn_w_mem[7358] = 68;
razn_w_mem[7359] = 68;
razn_w_mem[7360] = 68;
razn_w_mem[7361] = 68;
razn_w_mem[7362] = 68;
razn_w_mem[7363] = 68;
razn_w_mem[7364] = 68;
razn_w_mem[7365] = 68;
razn_w_mem[7366] = 68;
razn_w_mem[7367] = 68;
razn_w_mem[7368] = 68;
razn_w_mem[7369] = 68;
razn_w_mem[7370] = 68;
razn_w_mem[7371] = 68;
razn_w_mem[7372] = 68;
razn_w_mem[7373] = 68;
razn_w_mem[7374] = 68;
razn_w_mem[7375] = 68;
razn_w_mem[7376] = 68;
razn_w_mem[7377] = 68;
razn_w_mem[7378] = 68;
razn_w_mem[7379] = 68;
razn_w_mem[7380] = 68;
razn_w_mem[7381] = 68;
razn_w_mem[7382] = 68;
razn_w_mem[7383] = 68;
razn_w_mem[7384] = 68;
razn_w_mem[7385] = 68;
razn_w_mem[7386] = 68;
razn_w_mem[7387] = 68;
razn_w_mem[7388] = 68;
razn_w_mem[7389] = 68;
razn_w_mem[7390] = 68;
razn_w_mem[7391] = 68;
razn_w_mem[7392] = 68;
razn_w_mem[7393] = 68;
razn_w_mem[7394] = 68;
razn_w_mem[7395] = 68;
razn_w_mem[7396] = 68;
razn_w_mem[7397] = 68;
razn_w_mem[7398] = 68;
razn_w_mem[7399] = 68;
razn_w_mem[7400] = 68;
razn_w_mem[7401] = 68;
razn_w_mem[7402] = 68;
razn_w_mem[7403] = 68;
razn_w_mem[7404] = 68;
razn_w_mem[7405] = 68;
razn_w_mem[7406] = 68;
razn_w_mem[7407] = 68;
razn_w_mem[7408] = 68;
razn_w_mem[7409] = 68;
razn_w_mem[7410] = 68;
razn_w_mem[7411] = 68;
razn_w_mem[7412] = 68;
razn_w_mem[7413] = 68;
razn_w_mem[7414] = 68;
razn_w_mem[7415] = 68;
razn_w_mem[7416] = 68;
razn_w_mem[7417] = 68;
razn_w_mem[7418] = 68;
razn_w_mem[7419] = 68;
razn_w_mem[7420] = 68;
razn_w_mem[7421] = 68;
razn_w_mem[7422] = 68;
razn_w_mem[7423] = 68;
razn_w_mem[7424] = 38;
razn_w_mem[7425] = 38;
razn_w_mem[7426] = 38;
razn_w_mem[7427] = 38;
razn_w_mem[7428] = 38;
razn_w_mem[7429] = 38;
razn_w_mem[7430] = 38;
razn_w_mem[7431] = 38;
razn_w_mem[7432] = 38;
razn_w_mem[7433] = 38;
razn_w_mem[7434] = 38;
razn_w_mem[7435] = 38;
razn_w_mem[7436] = 38;
razn_w_mem[7437] = 38;
razn_w_mem[7438] = 38;
razn_w_mem[7439] = 38;
razn_w_mem[7440] = 38;
razn_w_mem[7441] = 38;
razn_w_mem[7442] = 38;
razn_w_mem[7443] = 38;
razn_w_mem[7444] = 38;
razn_w_mem[7445] = 38;
razn_w_mem[7446] = 38;
razn_w_mem[7447] = 38;
razn_w_mem[7448] = 38;
razn_w_mem[7449] = 38;
razn_w_mem[7450] = 38;
razn_w_mem[7451] = 38;
razn_w_mem[7452] = 38;
razn_w_mem[7453] = 38;
razn_w_mem[7454] = 38;
razn_w_mem[7455] = 38;
razn_w_mem[7456] = 38;
razn_w_mem[7457] = 38;
razn_w_mem[7458] = 38;
razn_w_mem[7459] = 38;
razn_w_mem[7460] = 38;
razn_w_mem[7461] = 38;
razn_w_mem[7462] = 38;
razn_w_mem[7463] = 38;
razn_w_mem[7464] = 38;
razn_w_mem[7465] = 38;
razn_w_mem[7466] = 38;
razn_w_mem[7467] = 38;
razn_w_mem[7468] = 38;
razn_w_mem[7469] = 38;
razn_w_mem[7470] = 38;
razn_w_mem[7471] = 38;
razn_w_mem[7472] = 38;
razn_w_mem[7473] = 38;
razn_w_mem[7474] = 38;
razn_w_mem[7475] = 38;
razn_w_mem[7476] = 38;
razn_w_mem[7477] = 38;
razn_w_mem[7478] = 38;
razn_w_mem[7479] = 38;
razn_w_mem[7480] = 38;
razn_w_mem[7481] = 38;
razn_w_mem[7482] = 38;
razn_w_mem[7483] = 38;
razn_w_mem[7484] = 38;
razn_w_mem[7485] = 38;
razn_w_mem[7486] = 38;
razn_w_mem[7487] = 38;
razn_w_mem[7488] = 38;
razn_w_mem[7489] = 38;
razn_w_mem[7490] = 38;
razn_w_mem[7491] = 38;
razn_w_mem[7492] = 38;
razn_w_mem[7493] = 38;
razn_w_mem[7494] = 38;
razn_w_mem[7495] = 38;
razn_w_mem[7496] = 38;
razn_w_mem[7497] = 38;
razn_w_mem[7498] = 38;
razn_w_mem[7499] = 38;
razn_w_mem[7500] = 38;
razn_w_mem[7501] = 38;
razn_w_mem[7502] = 38;
razn_w_mem[7503] = 38;
razn_w_mem[7504] = 38;
razn_w_mem[7505] = 38;
razn_w_mem[7506] = 38;
razn_w_mem[7507] = 38;
razn_w_mem[7508] = 38;
razn_w_mem[7509] = 38;
razn_w_mem[7510] = 38;
razn_w_mem[7511] = 38;
razn_w_mem[7512] = 38;
razn_w_mem[7513] = 38;
razn_w_mem[7514] = 38;
razn_w_mem[7515] = 38;
razn_w_mem[7516] = 38;
razn_w_mem[7517] = 38;
razn_w_mem[7518] = 38;
razn_w_mem[7519] = 38;
razn_w_mem[7520] = 38;
razn_w_mem[7521] = 38;
razn_w_mem[7522] = 38;
razn_w_mem[7523] = 38;
razn_w_mem[7524] = 38;
razn_w_mem[7525] = 38;
razn_w_mem[7526] = 38;
razn_w_mem[7527] = 38;
razn_w_mem[7528] = 38;
razn_w_mem[7529] = 38;
razn_w_mem[7530] = 38;
razn_w_mem[7531] = 38;
razn_w_mem[7532] = 38;
razn_w_mem[7533] = 38;
razn_w_mem[7534] = 38;
razn_w_mem[7535] = 38;
razn_w_mem[7536] = 38;
razn_w_mem[7537] = 38;
razn_w_mem[7538] = 38;
razn_w_mem[7539] = 38;
razn_w_mem[7540] = 38;
razn_w_mem[7541] = 38;
razn_w_mem[7542] = 38;
razn_w_mem[7543] = 38;
razn_w_mem[7544] = 38;
razn_w_mem[7545] = 38;
razn_w_mem[7546] = 38;
razn_w_mem[7547] = 38;
razn_w_mem[7548] = 38;
razn_w_mem[7549] = 38;
razn_w_mem[7550] = 38;
razn_w_mem[7551] = 38;
razn_w_mem[7552] = 8;
razn_w_mem[7553] = 8;
razn_w_mem[7554] = 8;
razn_w_mem[7555] = 8;
razn_w_mem[7556] = 8;
razn_w_mem[7557] = 8;
razn_w_mem[7558] = 8;
razn_w_mem[7559] = 8;
razn_w_mem[7560] = 8;
razn_w_mem[7561] = 8;
razn_w_mem[7562] = 8;
razn_w_mem[7563] = 8;
razn_w_mem[7564] = 8;
razn_w_mem[7565] = 8;
razn_w_mem[7566] = 8;
razn_w_mem[7567] = 8;
razn_w_mem[7568] = 8;
razn_w_mem[7569] = 8;
razn_w_mem[7570] = 8;
razn_w_mem[7571] = 8;
razn_w_mem[7572] = 8;
razn_w_mem[7573] = 8;
razn_w_mem[7574] = 8;
razn_w_mem[7575] = 8;
razn_w_mem[7576] = 8;
razn_w_mem[7577] = 8;
razn_w_mem[7578] = 8;
razn_w_mem[7579] = 8;
razn_w_mem[7580] = 8;
razn_w_mem[7581] = 8;
razn_w_mem[7582] = 8;
razn_w_mem[7583] = 8;
razn_w_mem[7584] = 8;
razn_w_mem[7585] = 8;
razn_w_mem[7586] = 8;
razn_w_mem[7587] = 8;
razn_w_mem[7588] = 8;
razn_w_mem[7589] = 8;
razn_w_mem[7590] = 8;
razn_w_mem[7591] = 8;
razn_w_mem[7592] = 8;
razn_w_mem[7593] = 8;
razn_w_mem[7594] = 8;
razn_w_mem[7595] = 8;
razn_w_mem[7596] = 8;
razn_w_mem[7597] = 8;
razn_w_mem[7598] = 8;
razn_w_mem[7599] = 8;
razn_w_mem[7600] = 8;
razn_w_mem[7601] = 8;
razn_w_mem[7602] = 8;
razn_w_mem[7603] = 8;
razn_w_mem[7604] = 8;
razn_w_mem[7605] = 8;
razn_w_mem[7606] = 8;
razn_w_mem[7607] = 8;
razn_w_mem[7608] = 8;
razn_w_mem[7609] = 8;
razn_w_mem[7610] = 8;
razn_w_mem[7611] = 8;
razn_w_mem[7612] = 8;
razn_w_mem[7613] = 8;
razn_w_mem[7614] = 8;
razn_w_mem[7615] = 8;
razn_w_mem[7616] = 8;
razn_w_mem[7617] = 8;
razn_w_mem[7618] = 8;
razn_w_mem[7619] = 8;
razn_w_mem[7620] = 8;
razn_w_mem[7621] = 8;
razn_w_mem[7622] = 8;
razn_w_mem[7623] = 8;
razn_w_mem[7624] = 8;
razn_w_mem[7625] = 8;
razn_w_mem[7626] = 8;
razn_w_mem[7627] = 8;
razn_w_mem[7628] = 8;
razn_w_mem[7629] = 8;
razn_w_mem[7630] = 8;
razn_w_mem[7631] = 8;
razn_w_mem[7632] = 8;
razn_w_mem[7633] = 8;
razn_w_mem[7634] = 8;
razn_w_mem[7635] = 8;
razn_w_mem[7636] = 8;
razn_w_mem[7637] = 8;
razn_w_mem[7638] = 8;
razn_w_mem[7639] = 8;
razn_w_mem[7640] = 8;
razn_w_mem[7641] = 8;
razn_w_mem[7642] = 8;
razn_w_mem[7643] = 8;
razn_w_mem[7644] = 8;
razn_w_mem[7645] = 8;
razn_w_mem[7646] = 8;
razn_w_mem[7647] = 8;
razn_w_mem[7648] = 8;
razn_w_mem[7649] = 8;
razn_w_mem[7650] = 8;
razn_w_mem[7651] = 8;
razn_w_mem[7652] = 8;
razn_w_mem[7653] = 8;
razn_w_mem[7654] = 8;
razn_w_mem[7655] = 8;
razn_w_mem[7656] = 8;
razn_w_mem[7657] = 8;
razn_w_mem[7658] = 8;
razn_w_mem[7659] = 8;
razn_w_mem[7660] = 8;
razn_w_mem[7661] = 8;
razn_w_mem[7662] = 8;
razn_w_mem[7663] = 8;
razn_w_mem[7664] = 8;
razn_w_mem[7665] = 8;
razn_w_mem[7666] = 8;
razn_w_mem[7667] = 8;
razn_w_mem[7668] = 8;
razn_w_mem[7669] = 8;
razn_w_mem[7670] = 8;
razn_w_mem[7671] = 8;
razn_w_mem[7672] = 8;
razn_w_mem[7673] = 8;
razn_w_mem[7674] = 8;
razn_w_mem[7675] = 8;
razn_w_mem[7676] = 8;
razn_w_mem[7677] = 8;
razn_w_mem[7678] = 8;
razn_w_mem[7679] = 8;
razn_w_mem[7680] = 232;
razn_w_mem[7681] = 232;
razn_w_mem[7682] = 232;
razn_w_mem[7683] = 232;
razn_w_mem[7684] = 232;
razn_w_mem[7685] = 232;
razn_w_mem[7686] = 232;
razn_w_mem[7687] = 232;
razn_w_mem[7688] = 232;
razn_w_mem[7689] = 232;
razn_w_mem[7690] = 232;
razn_w_mem[7691] = 232;
razn_w_mem[7692] = 232;
razn_w_mem[7693] = 232;
razn_w_mem[7694] = 232;
razn_w_mem[7695] = 232;
razn_w_mem[7696] = 232;
razn_w_mem[7697] = 232;
razn_w_mem[7698] = 232;
razn_w_mem[7699] = 232;
razn_w_mem[7700] = 232;
razn_w_mem[7701] = 232;
razn_w_mem[7702] = 232;
razn_w_mem[7703] = 232;
razn_w_mem[7704] = 232;
razn_w_mem[7705] = 232;
razn_w_mem[7706] = 232;
razn_w_mem[7707] = 232;
razn_w_mem[7708] = 232;
razn_w_mem[7709] = 232;
razn_w_mem[7710] = 232;
razn_w_mem[7711] = 232;
razn_w_mem[7712] = 232;
razn_w_mem[7713] = 232;
razn_w_mem[7714] = 232;
razn_w_mem[7715] = 232;
razn_w_mem[7716] = 232;
razn_w_mem[7717] = 232;
razn_w_mem[7718] = 232;
razn_w_mem[7719] = 232;
razn_w_mem[7720] = 232;
razn_w_mem[7721] = 232;
razn_w_mem[7722] = 232;
razn_w_mem[7723] = 232;
razn_w_mem[7724] = 232;
razn_w_mem[7725] = 232;
razn_w_mem[7726] = 232;
razn_w_mem[7727] = 232;
razn_w_mem[7728] = 232;
razn_w_mem[7729] = 232;
razn_w_mem[7730] = 232;
razn_w_mem[7731] = 232;
razn_w_mem[7732] = 232;
razn_w_mem[7733] = 232;
razn_w_mem[7734] = 232;
razn_w_mem[7735] = 232;
razn_w_mem[7736] = 232;
razn_w_mem[7737] = 232;
razn_w_mem[7738] = 232;
razn_w_mem[7739] = 232;
razn_w_mem[7740] = 232;
razn_w_mem[7741] = 232;
razn_w_mem[7742] = 232;
razn_w_mem[7743] = 232;
razn_w_mem[7744] = 232;
razn_w_mem[7745] = 232;
razn_w_mem[7746] = 232;
razn_w_mem[7747] = 232;
razn_w_mem[7748] = 232;
razn_w_mem[7749] = 232;
razn_w_mem[7750] = 232;
razn_w_mem[7751] = 232;
razn_w_mem[7752] = 232;
razn_w_mem[7753] = 232;
razn_w_mem[7754] = 232;
razn_w_mem[7755] = 232;
razn_w_mem[7756] = 232;
razn_w_mem[7757] = 232;
razn_w_mem[7758] = 232;
razn_w_mem[7759] = 232;
razn_w_mem[7760] = 232;
razn_w_mem[7761] = 232;
razn_w_mem[7762] = 232;
razn_w_mem[7763] = 232;
razn_w_mem[7764] = 232;
razn_w_mem[7765] = 232;
razn_w_mem[7766] = 232;
razn_w_mem[7767] = 232;
razn_w_mem[7768] = 232;
razn_w_mem[7769] = 232;
razn_w_mem[7770] = 232;
razn_w_mem[7771] = 232;
razn_w_mem[7772] = 232;
razn_w_mem[7773] = 232;
razn_w_mem[7774] = 232;
razn_w_mem[7775] = 232;
razn_w_mem[7776] = 232;
razn_w_mem[7777] = 232;
razn_w_mem[7778] = 232;
razn_w_mem[7779] = 232;
razn_w_mem[7780] = 232;
razn_w_mem[7781] = 232;
razn_w_mem[7782] = 232;
razn_w_mem[7783] = 232;
razn_w_mem[7784] = 232;
razn_w_mem[7785] = 232;
razn_w_mem[7786] = 232;
razn_w_mem[7787] = 232;
razn_w_mem[7788] = 232;
razn_w_mem[7789] = 232;
razn_w_mem[7790] = 232;
razn_w_mem[7791] = 232;
razn_w_mem[7792] = 232;
razn_w_mem[7793] = 232;
razn_w_mem[7794] = 232;
razn_w_mem[7795] = 232;
razn_w_mem[7796] = 232;
razn_w_mem[7797] = 232;
razn_w_mem[7798] = 232;
razn_w_mem[7799] = 232;
razn_w_mem[7800] = 232;
razn_w_mem[7801] = 232;
razn_w_mem[7802] = 232;
razn_w_mem[7803] = 232;
razn_w_mem[7804] = 232;
razn_w_mem[7805] = 232;
razn_w_mem[7806] = 232;
razn_w_mem[7807] = 232;
razn_w_mem[7808] = 202;
razn_w_mem[7809] = 202;
razn_w_mem[7810] = 202;
razn_w_mem[7811] = 202;
razn_w_mem[7812] = 202;
razn_w_mem[7813] = 202;
razn_w_mem[7814] = 202;
razn_w_mem[7815] = 202;
razn_w_mem[7816] = 202;
razn_w_mem[7817] = 202;
razn_w_mem[7818] = 202;
razn_w_mem[7819] = 202;
razn_w_mem[7820] = 202;
razn_w_mem[7821] = 202;
razn_w_mem[7822] = 202;
razn_w_mem[7823] = 202;
razn_w_mem[7824] = 202;
razn_w_mem[7825] = 202;
razn_w_mem[7826] = 202;
razn_w_mem[7827] = 202;
razn_w_mem[7828] = 202;
razn_w_mem[7829] = 202;
razn_w_mem[7830] = 202;
razn_w_mem[7831] = 202;
razn_w_mem[7832] = 202;
razn_w_mem[7833] = 202;
razn_w_mem[7834] = 202;
razn_w_mem[7835] = 202;
razn_w_mem[7836] = 202;
razn_w_mem[7837] = 202;
razn_w_mem[7838] = 202;
razn_w_mem[7839] = 202;
razn_w_mem[7840] = 202;
razn_w_mem[7841] = 202;
razn_w_mem[7842] = 202;
razn_w_mem[7843] = 202;
razn_w_mem[7844] = 202;
razn_w_mem[7845] = 202;
razn_w_mem[7846] = 202;
razn_w_mem[7847] = 202;
razn_w_mem[7848] = 202;
razn_w_mem[7849] = 202;
razn_w_mem[7850] = 202;
razn_w_mem[7851] = 202;
razn_w_mem[7852] = 202;
razn_w_mem[7853] = 202;
razn_w_mem[7854] = 202;
razn_w_mem[7855] = 202;
razn_w_mem[7856] = 202;
razn_w_mem[7857] = 202;
razn_w_mem[7858] = 202;
razn_w_mem[7859] = 202;
razn_w_mem[7860] = 202;
razn_w_mem[7861] = 202;
razn_w_mem[7862] = 202;
razn_w_mem[7863] = 202;
razn_w_mem[7864] = 202;
razn_w_mem[7865] = 202;
razn_w_mem[7866] = 202;
razn_w_mem[7867] = 202;
razn_w_mem[7868] = 202;
razn_w_mem[7869] = 202;
razn_w_mem[7870] = 202;
razn_w_mem[7871] = 202;
razn_w_mem[7872] = 202;
razn_w_mem[7873] = 202;
razn_w_mem[7874] = 202;
razn_w_mem[7875] = 202;
razn_w_mem[7876] = 202;
razn_w_mem[7877] = 202;
razn_w_mem[7878] = 202;
razn_w_mem[7879] = 202;
razn_w_mem[7880] = 202;
razn_w_mem[7881] = 202;
razn_w_mem[7882] = 202;
razn_w_mem[7883] = 202;
razn_w_mem[7884] = 202;
razn_w_mem[7885] = 202;
razn_w_mem[7886] = 202;
razn_w_mem[7887] = 202;
razn_w_mem[7888] = 202;
razn_w_mem[7889] = 202;
razn_w_mem[7890] = 202;
razn_w_mem[7891] = 202;
razn_w_mem[7892] = 202;
razn_w_mem[7893] = 202;
razn_w_mem[7894] = 202;
razn_w_mem[7895] = 202;
razn_w_mem[7896] = 202;
razn_w_mem[7897] = 202;
razn_w_mem[7898] = 202;
razn_w_mem[7899] = 202;
razn_w_mem[7900] = 202;
razn_w_mem[7901] = 202;
razn_w_mem[7902] = 202;
razn_w_mem[7903] = 202;
razn_w_mem[7904] = 202;
razn_w_mem[7905] = 202;
razn_w_mem[7906] = 202;
razn_w_mem[7907] = 202;
razn_w_mem[7908] = 202;
razn_w_mem[7909] = 202;
razn_w_mem[7910] = 202;
razn_w_mem[7911] = 202;
razn_w_mem[7912] = 202;
razn_w_mem[7913] = 202;
razn_w_mem[7914] = 202;
razn_w_mem[7915] = 202;
razn_w_mem[7916] = 202;
razn_w_mem[7917] = 202;
razn_w_mem[7918] = 202;
razn_w_mem[7919] = 202;
razn_w_mem[7920] = 202;
razn_w_mem[7921] = 202;
razn_w_mem[7922] = 202;
razn_w_mem[7923] = 202;
razn_w_mem[7924] = 202;
razn_w_mem[7925] = 202;
razn_w_mem[7926] = 202;
razn_w_mem[7927] = 202;
razn_w_mem[7928] = 202;
razn_w_mem[7929] = 202;
razn_w_mem[7930] = 202;
razn_w_mem[7931] = 202;
razn_w_mem[7932] = 202;
razn_w_mem[7933] = 202;
razn_w_mem[7934] = 202;
razn_w_mem[7935] = 202;
razn_w_mem[7936] = 172;
razn_w_mem[7937] = 172;
razn_w_mem[7938] = 172;
razn_w_mem[7939] = 172;
razn_w_mem[7940] = 172;
razn_w_mem[7941] = 172;
razn_w_mem[7942] = 172;
razn_w_mem[7943] = 172;
razn_w_mem[7944] = 172;
razn_w_mem[7945] = 172;
razn_w_mem[7946] = 172;
razn_w_mem[7947] = 172;
razn_w_mem[7948] = 172;
razn_w_mem[7949] = 172;
razn_w_mem[7950] = 172;
razn_w_mem[7951] = 172;
razn_w_mem[7952] = 172;
razn_w_mem[7953] = 172;
razn_w_mem[7954] = 172;
razn_w_mem[7955] = 172;
razn_w_mem[7956] = 172;
razn_w_mem[7957] = 172;
razn_w_mem[7958] = 172;
razn_w_mem[7959] = 172;
razn_w_mem[7960] = 172;
razn_w_mem[7961] = 172;
razn_w_mem[7962] = 172;
razn_w_mem[7963] = 172;
razn_w_mem[7964] = 172;
razn_w_mem[7965] = 172;
razn_w_mem[7966] = 172;
razn_w_mem[7967] = 172;
razn_w_mem[7968] = 172;
razn_w_mem[7969] = 172;
razn_w_mem[7970] = 172;
razn_w_mem[7971] = 172;
razn_w_mem[7972] = 172;
razn_w_mem[7973] = 172;
razn_w_mem[7974] = 172;
razn_w_mem[7975] = 172;
razn_w_mem[7976] = 172;
razn_w_mem[7977] = 172;
razn_w_mem[7978] = 172;
razn_w_mem[7979] = 172;
razn_w_mem[7980] = 172;
razn_w_mem[7981] = 172;
razn_w_mem[7982] = 172;
razn_w_mem[7983] = 172;
razn_w_mem[7984] = 172;
razn_w_mem[7985] = 172;
razn_w_mem[7986] = 172;
razn_w_mem[7987] = 172;
razn_w_mem[7988] = 172;
razn_w_mem[7989] = 172;
razn_w_mem[7990] = 172;
razn_w_mem[7991] = 172;
razn_w_mem[7992] = 172;
razn_w_mem[7993] = 172;
razn_w_mem[7994] = 172;
razn_w_mem[7995] = 172;
razn_w_mem[7996] = 172;
razn_w_mem[7997] = 172;
razn_w_mem[7998] = 172;
razn_w_mem[7999] = 172;
razn_w_mem[8000] = 172;
razn_w_mem[8001] = 172;
razn_w_mem[8002] = 172;
razn_w_mem[8003] = 172;
razn_w_mem[8004] = 172;
razn_w_mem[8005] = 172;
razn_w_mem[8006] = 172;
razn_w_mem[8007] = 172;
razn_w_mem[8008] = 172;
razn_w_mem[8009] = 172;
razn_w_mem[8010] = 172;
razn_w_mem[8011] = 172;
razn_w_mem[8012] = 172;
razn_w_mem[8013] = 172;
razn_w_mem[8014] = 172;
razn_w_mem[8015] = 172;
razn_w_mem[8016] = 172;
razn_w_mem[8017] = 172;
razn_w_mem[8018] = 172;
razn_w_mem[8019] = 172;
razn_w_mem[8020] = 172;
razn_w_mem[8021] = 172;
razn_w_mem[8022] = 172;
razn_w_mem[8023] = 172;
razn_w_mem[8024] = 172;
razn_w_mem[8025] = 172;
razn_w_mem[8026] = 172;
razn_w_mem[8027] = 172;
razn_w_mem[8028] = 172;
razn_w_mem[8029] = 172;
razn_w_mem[8030] = 172;
razn_w_mem[8031] = 172;
razn_w_mem[8032] = 172;
razn_w_mem[8033] = 172;
razn_w_mem[8034] = 172;
razn_w_mem[8035] = 172;
razn_w_mem[8036] = 172;
razn_w_mem[8037] = 172;
razn_w_mem[8038] = 172;
razn_w_mem[8039] = 172;
razn_w_mem[8040] = 172;
razn_w_mem[8041] = 172;
razn_w_mem[8042] = 172;
razn_w_mem[8043] = 172;
razn_w_mem[8044] = 172;
razn_w_mem[8045] = 172;
razn_w_mem[8046] = 172;
razn_w_mem[8047] = 172;
razn_w_mem[8048] = 172;
razn_w_mem[8049] = 172;
razn_w_mem[8050] = 172;
razn_w_mem[8051] = 172;
razn_w_mem[8052] = 172;
razn_w_mem[8053] = 172;
razn_w_mem[8054] = 172;
razn_w_mem[8055] = 172;
razn_w_mem[8056] = 172;
razn_w_mem[8057] = 172;
razn_w_mem[8058] = 172;
razn_w_mem[8059] = 172;
razn_w_mem[8060] = 172;
razn_w_mem[8061] = 172;
razn_w_mem[8062] = 172;
razn_w_mem[8063] = 172;
razn_w_mem[8064] = 142;
razn_w_mem[8065] = 142;
razn_w_mem[8066] = 142;
razn_w_mem[8067] = 142;
razn_w_mem[8068] = 142;
razn_w_mem[8069] = 142;
razn_w_mem[8070] = 142;
razn_w_mem[8071] = 142;
razn_w_mem[8072] = 142;
razn_w_mem[8073] = 142;
razn_w_mem[8074] = 142;
razn_w_mem[8075] = 142;
razn_w_mem[8076] = 142;
razn_w_mem[8077] = 142;
razn_w_mem[8078] = 142;
razn_w_mem[8079] = 142;
razn_w_mem[8080] = 142;
razn_w_mem[8081] = 142;
razn_w_mem[8082] = 142;
razn_w_mem[8083] = 142;
razn_w_mem[8084] = 142;
razn_w_mem[8085] = 142;
razn_w_mem[8086] = 142;
razn_w_mem[8087] = 142;
razn_w_mem[8088] = 142;
razn_w_mem[8089] = 142;
razn_w_mem[8090] = 142;
razn_w_mem[8091] = 142;
razn_w_mem[8092] = 142;
razn_w_mem[8093] = 142;
razn_w_mem[8094] = 142;
razn_w_mem[8095] = 142;
razn_w_mem[8096] = 142;
razn_w_mem[8097] = 142;
razn_w_mem[8098] = 142;
razn_w_mem[8099] = 142;
razn_w_mem[8100] = 142;
razn_w_mem[8101] = 142;
razn_w_mem[8102] = 142;
razn_w_mem[8103] = 142;
razn_w_mem[8104] = 142;
razn_w_mem[8105] = 142;
razn_w_mem[8106] = 142;
razn_w_mem[8107] = 142;
razn_w_mem[8108] = 142;
razn_w_mem[8109] = 142;
razn_w_mem[8110] = 142;
razn_w_mem[8111] = 142;
razn_w_mem[8112] = 142;
razn_w_mem[8113] = 142;
razn_w_mem[8114] = 142;
razn_w_mem[8115] = 142;
razn_w_mem[8116] = 142;
razn_w_mem[8117] = 142;
razn_w_mem[8118] = 142;
razn_w_mem[8119] = 142;
razn_w_mem[8120] = 142;
razn_w_mem[8121] = 142;
razn_w_mem[8122] = 142;
razn_w_mem[8123] = 142;
razn_w_mem[8124] = 142;
razn_w_mem[8125] = 142;
razn_w_mem[8126] = 142;
razn_w_mem[8127] = 142;
razn_w_mem[8128] = 142;
razn_w_mem[8129] = 142;
razn_w_mem[8130] = 142;
razn_w_mem[8131] = 142;
razn_w_mem[8132] = 142;
razn_w_mem[8133] = 142;
razn_w_mem[8134] = 142;
razn_w_mem[8135] = 142;
razn_w_mem[8136] = 142;
razn_w_mem[8137] = 142;
razn_w_mem[8138] = 142;
razn_w_mem[8139] = 142;
razn_w_mem[8140] = 142;
razn_w_mem[8141] = 142;
razn_w_mem[8142] = 142;
razn_w_mem[8143] = 142;
razn_w_mem[8144] = 142;
razn_w_mem[8145] = 142;
razn_w_mem[8146] = 142;
razn_w_mem[8147] = 142;
razn_w_mem[8148] = 142;
razn_w_mem[8149] = 142;
razn_w_mem[8150] = 142;
razn_w_mem[8151] = 142;
razn_w_mem[8152] = 142;
razn_w_mem[8153] = 142;
razn_w_mem[8154] = 142;
razn_w_mem[8155] = 142;
razn_w_mem[8156] = 142;
razn_w_mem[8157] = 142;
razn_w_mem[8158] = 142;
razn_w_mem[8159] = 142;
razn_w_mem[8160] = 142;
razn_w_mem[8161] = 142;
razn_w_mem[8162] = 142;
razn_w_mem[8163] = 142;
razn_w_mem[8164] = 142;
razn_w_mem[8165] = 142;
razn_w_mem[8166] = 142;
razn_w_mem[8167] = 142;
razn_w_mem[8168] = 142;
razn_w_mem[8169] = 142;
razn_w_mem[8170] = 142;
razn_w_mem[8171] = 142;
razn_w_mem[8172] = 142;
razn_w_mem[8173] = 142;
razn_w_mem[8174] = 142;
razn_w_mem[8175] = 142;
razn_w_mem[8176] = 142;
razn_w_mem[8177] = 142;
razn_w_mem[8178] = 142;
razn_w_mem[8179] = 142;
razn_w_mem[8180] = 142;
razn_w_mem[8181] = 142;
razn_w_mem[8182] = 142;
razn_w_mem[8183] = 142;
razn_w_mem[8184] = 142;
razn_w_mem[8185] = 142;
razn_w_mem[8186] = 142;
razn_w_mem[8187] = 142;
razn_w_mem[8188] = 142;
razn_w_mem[8189] = 142;
razn_w_mem[8190] = 142;
razn_w_mem[8191] = 142;
razn_w_mem[8192] = 112;
razn_w_mem[8193] = 112;
razn_w_mem[8194] = 112;
razn_w_mem[8195] = 112;
razn_w_mem[8196] = 112;
razn_w_mem[8197] = 112;
razn_w_mem[8198] = 112;
razn_w_mem[8199] = 112;
razn_w_mem[8200] = 112;
razn_w_mem[8201] = 112;
razn_w_mem[8202] = 112;
razn_w_mem[8203] = 112;
razn_w_mem[8204] = 112;
razn_w_mem[8205] = 112;
razn_w_mem[8206] = 112;
razn_w_mem[8207] = 112;
razn_w_mem[8208] = 112;
razn_w_mem[8209] = 112;
razn_w_mem[8210] = 112;
razn_w_mem[8211] = 112;
razn_w_mem[8212] = 112;
razn_w_mem[8213] = 112;
razn_w_mem[8214] = 112;
razn_w_mem[8215] = 112;
razn_w_mem[8216] = 112;
razn_w_mem[8217] = 112;
razn_w_mem[8218] = 112;
razn_w_mem[8219] = 112;
razn_w_mem[8220] = 112;
razn_w_mem[8221] = 112;
razn_w_mem[8222] = 112;
razn_w_mem[8223] = 112;
razn_w_mem[8224] = 112;
razn_w_mem[8225] = 112;
razn_w_mem[8226] = 112;
razn_w_mem[8227] = 112;
razn_w_mem[8228] = 112;
razn_w_mem[8229] = 112;
razn_w_mem[8230] = 112;
razn_w_mem[8231] = 112;
razn_w_mem[8232] = 112;
razn_w_mem[8233] = 112;
razn_w_mem[8234] = 112;
razn_w_mem[8235] = 112;
razn_w_mem[8236] = 112;
razn_w_mem[8237] = 112;
razn_w_mem[8238] = 112;
razn_w_mem[8239] = 112;
razn_w_mem[8240] = 112;
razn_w_mem[8241] = 112;
razn_w_mem[8242] = 112;
razn_w_mem[8243] = 112;
razn_w_mem[8244] = 112;
razn_w_mem[8245] = 112;
razn_w_mem[8246] = 112;
razn_w_mem[8247] = 112;
razn_w_mem[8248] = 112;
razn_w_mem[8249] = 112;
razn_w_mem[8250] = 112;
razn_w_mem[8251] = 112;
razn_w_mem[8252] = 112;
razn_w_mem[8253] = 112;
razn_w_mem[8254] = 112;
razn_w_mem[8255] = 112;
razn_w_mem[8256] = 112;
razn_w_mem[8257] = 112;
razn_w_mem[8258] = 112;
razn_w_mem[8259] = 112;
razn_w_mem[8260] = 112;
razn_w_mem[8261] = 112;
razn_w_mem[8262] = 112;
razn_w_mem[8263] = 112;
razn_w_mem[8264] = 112;
razn_w_mem[8265] = 112;
razn_w_mem[8266] = 112;
razn_w_mem[8267] = 112;
razn_w_mem[8268] = 112;
razn_w_mem[8269] = 112;
razn_w_mem[8270] = 112;
razn_w_mem[8271] = 112;
razn_w_mem[8272] = 112;
razn_w_mem[8273] = 112;
razn_w_mem[8274] = 112;
razn_w_mem[8275] = 112;
razn_w_mem[8276] = 112;
razn_w_mem[8277] = 112;
razn_w_mem[8278] = 112;
razn_w_mem[8279] = 112;
razn_w_mem[8280] = 112;
razn_w_mem[8281] = 112;
razn_w_mem[8282] = 112;
razn_w_mem[8283] = 112;
razn_w_mem[8284] = 112;
razn_w_mem[8285] = 112;
razn_w_mem[8286] = 112;
razn_w_mem[8287] = 112;
razn_w_mem[8288] = 112;
razn_w_mem[8289] = 112;
razn_w_mem[8290] = 112;
razn_w_mem[8291] = 112;
razn_w_mem[8292] = 112;
razn_w_mem[8293] = 112;
razn_w_mem[8294] = 112;
razn_w_mem[8295] = 112;
razn_w_mem[8296] = 112;
razn_w_mem[8297] = 112;
razn_w_mem[8298] = 112;
razn_w_mem[8299] = 112;
razn_w_mem[8300] = 112;
razn_w_mem[8301] = 112;
razn_w_mem[8302] = 112;
razn_w_mem[8303] = 112;
razn_w_mem[8304] = 112;
razn_w_mem[8305] = 112;
razn_w_mem[8306] = 112;
razn_w_mem[8307] = 112;
razn_w_mem[8308] = 112;
razn_w_mem[8309] = 112;
razn_w_mem[8310] = 112;
razn_w_mem[8311] = 112;
razn_w_mem[8312] = 112;
razn_w_mem[8313] = 112;
razn_w_mem[8314] = 112;
razn_w_mem[8315] = 112;
razn_w_mem[8316] = 112;
razn_w_mem[8317] = 112;
razn_w_mem[8318] = 112;
razn_w_mem[8319] = 112;
razn_w_mem[8320] = 82;
razn_w_mem[8321] = 82;
razn_w_mem[8322] = 82;
razn_w_mem[8323] = 82;
razn_w_mem[8324] = 82;
razn_w_mem[8325] = 82;
razn_w_mem[8326] = 82;
razn_w_mem[8327] = 82;
razn_w_mem[8328] = 82;
razn_w_mem[8329] = 82;
razn_w_mem[8330] = 82;
razn_w_mem[8331] = 82;
razn_w_mem[8332] = 82;
razn_w_mem[8333] = 82;
razn_w_mem[8334] = 82;
razn_w_mem[8335] = 82;
razn_w_mem[8336] = 82;
razn_w_mem[8337] = 82;
razn_w_mem[8338] = 82;
razn_w_mem[8339] = 82;
razn_w_mem[8340] = 82;
razn_w_mem[8341] = 82;
razn_w_mem[8342] = 82;
razn_w_mem[8343] = 82;
razn_w_mem[8344] = 82;
razn_w_mem[8345] = 82;
razn_w_mem[8346] = 82;
razn_w_mem[8347] = 82;
razn_w_mem[8348] = 82;
razn_w_mem[8349] = 82;
razn_w_mem[8350] = 82;
razn_w_mem[8351] = 82;
razn_w_mem[8352] = 82;
razn_w_mem[8353] = 82;
razn_w_mem[8354] = 82;
razn_w_mem[8355] = 82;
razn_w_mem[8356] = 82;
razn_w_mem[8357] = 82;
razn_w_mem[8358] = 82;
razn_w_mem[8359] = 82;
razn_w_mem[8360] = 82;
razn_w_mem[8361] = 82;
razn_w_mem[8362] = 82;
razn_w_mem[8363] = 82;
razn_w_mem[8364] = 82;
razn_w_mem[8365] = 82;
razn_w_mem[8366] = 82;
razn_w_mem[8367] = 82;
razn_w_mem[8368] = 82;
razn_w_mem[8369] = 82;
razn_w_mem[8370] = 82;
razn_w_mem[8371] = 82;
razn_w_mem[8372] = 82;
razn_w_mem[8373] = 82;
razn_w_mem[8374] = 82;
razn_w_mem[8375] = 82;
razn_w_mem[8376] = 82;
razn_w_mem[8377] = 82;
razn_w_mem[8378] = 82;
razn_w_mem[8379] = 82;
razn_w_mem[8380] = 82;
razn_w_mem[8381] = 82;
razn_w_mem[8382] = 82;
razn_w_mem[8383] = 82;
razn_w_mem[8384] = 82;
razn_w_mem[8385] = 82;
razn_w_mem[8386] = 82;
razn_w_mem[8387] = 82;
razn_w_mem[8388] = 82;
razn_w_mem[8389] = 82;
razn_w_mem[8390] = 82;
razn_w_mem[8391] = 82;
razn_w_mem[8392] = 82;
razn_w_mem[8393] = 82;
razn_w_mem[8394] = 82;
razn_w_mem[8395] = 82;
razn_w_mem[8396] = 82;
razn_w_mem[8397] = 82;
razn_w_mem[8398] = 82;
razn_w_mem[8399] = 82;
razn_w_mem[8400] = 82;
razn_w_mem[8401] = 82;
razn_w_mem[8402] = 82;
razn_w_mem[8403] = 82;
razn_w_mem[8404] = 82;
razn_w_mem[8405] = 82;
razn_w_mem[8406] = 82;
razn_w_mem[8407] = 82;
razn_w_mem[8408] = 82;
razn_w_mem[8409] = 82;
razn_w_mem[8410] = 82;
razn_w_mem[8411] = 82;
razn_w_mem[8412] = 82;
razn_w_mem[8413] = 82;
razn_w_mem[8414] = 82;
razn_w_mem[8415] = 82;
razn_w_mem[8416] = 82;
razn_w_mem[8417] = 82;
razn_w_mem[8418] = 82;
razn_w_mem[8419] = 82;
razn_w_mem[8420] = 82;
razn_w_mem[8421] = 82;
razn_w_mem[8422] = 82;
razn_w_mem[8423] = 82;
razn_w_mem[8424] = 82;
razn_w_mem[8425] = 82;
razn_w_mem[8426] = 82;
razn_w_mem[8427] = 82;
razn_w_mem[8428] = 82;
razn_w_mem[8429] = 82;
razn_w_mem[8430] = 82;
razn_w_mem[8431] = 82;
razn_w_mem[8432] = 82;
razn_w_mem[8433] = 82;
razn_w_mem[8434] = 82;
razn_w_mem[8435] = 82;
razn_w_mem[8436] = 82;
razn_w_mem[8437] = 82;
razn_w_mem[8438] = 82;
razn_w_mem[8439] = 82;
razn_w_mem[8440] = 82;
razn_w_mem[8441] = 82;
razn_w_mem[8442] = 82;
razn_w_mem[8443] = 82;
razn_w_mem[8444] = 82;
razn_w_mem[8445] = 82;
razn_w_mem[8446] = 82;
razn_w_mem[8447] = 82;
razn_w_mem[8448] = 52;
razn_w_mem[8449] = 52;
razn_w_mem[8450] = 52;
razn_w_mem[8451] = 52;
razn_w_mem[8452] = 52;
razn_w_mem[8453] = 52;
razn_w_mem[8454] = 52;
razn_w_mem[8455] = 52;
razn_w_mem[8456] = 52;
razn_w_mem[8457] = 52;
razn_w_mem[8458] = 52;
razn_w_mem[8459] = 52;
razn_w_mem[8460] = 52;
razn_w_mem[8461] = 52;
razn_w_mem[8462] = 52;
razn_w_mem[8463] = 52;
razn_w_mem[8464] = 52;
razn_w_mem[8465] = 52;
razn_w_mem[8466] = 52;
razn_w_mem[8467] = 52;
razn_w_mem[8468] = 52;
razn_w_mem[8469] = 52;
razn_w_mem[8470] = 52;
razn_w_mem[8471] = 52;
razn_w_mem[8472] = 52;
razn_w_mem[8473] = 52;
razn_w_mem[8474] = 52;
razn_w_mem[8475] = 52;
razn_w_mem[8476] = 52;
razn_w_mem[8477] = 52;
razn_w_mem[8478] = 52;
razn_w_mem[8479] = 52;
razn_w_mem[8480] = 52;
razn_w_mem[8481] = 52;
razn_w_mem[8482] = 52;
razn_w_mem[8483] = 52;
razn_w_mem[8484] = 52;
razn_w_mem[8485] = 52;
razn_w_mem[8486] = 52;
razn_w_mem[8487] = 52;
razn_w_mem[8488] = 52;
razn_w_mem[8489] = 52;
razn_w_mem[8490] = 52;
razn_w_mem[8491] = 52;
razn_w_mem[8492] = 52;
razn_w_mem[8493] = 52;
razn_w_mem[8494] = 52;
razn_w_mem[8495] = 52;
razn_w_mem[8496] = 52;
razn_w_mem[8497] = 52;
razn_w_mem[8498] = 52;
razn_w_mem[8499] = 52;
razn_w_mem[8500] = 52;
razn_w_mem[8501] = 52;
razn_w_mem[8502] = 52;
razn_w_mem[8503] = 52;
razn_w_mem[8504] = 52;
razn_w_mem[8505] = 52;
razn_w_mem[8506] = 52;
razn_w_mem[8507] = 52;
razn_w_mem[8508] = 52;
razn_w_mem[8509] = 52;
razn_w_mem[8510] = 52;
razn_w_mem[8511] = 52;
razn_w_mem[8512] = 52;
razn_w_mem[8513] = 52;
razn_w_mem[8514] = 52;
razn_w_mem[8515] = 52;
razn_w_mem[8516] = 52;
razn_w_mem[8517] = 52;
razn_w_mem[8518] = 52;
razn_w_mem[8519] = 52;
razn_w_mem[8520] = 52;
razn_w_mem[8521] = 52;
razn_w_mem[8522] = 52;
razn_w_mem[8523] = 52;
razn_w_mem[8524] = 52;
razn_w_mem[8525] = 52;
razn_w_mem[8526] = 52;
razn_w_mem[8527] = 52;
razn_w_mem[8528] = 52;
razn_w_mem[8529] = 52;
razn_w_mem[8530] = 52;
razn_w_mem[8531] = 52;
razn_w_mem[8532] = 52;
razn_w_mem[8533] = 52;
razn_w_mem[8534] = 52;
razn_w_mem[8535] = 52;
razn_w_mem[8536] = 52;
razn_w_mem[8537] = 52;
razn_w_mem[8538] = 52;
razn_w_mem[8539] = 52;
razn_w_mem[8540] = 52;
razn_w_mem[8541] = 52;
razn_w_mem[8542] = 52;
razn_w_mem[8543] = 52;
razn_w_mem[8544] = 52;
razn_w_mem[8545] = 52;
razn_w_mem[8546] = 52;
razn_w_mem[8547] = 52;
razn_w_mem[8548] = 52;
razn_w_mem[8549] = 52;
razn_w_mem[8550] = 52;
razn_w_mem[8551] = 52;
razn_w_mem[8552] = 52;
razn_w_mem[8553] = 52;
razn_w_mem[8554] = 52;
razn_w_mem[8555] = 52;
razn_w_mem[8556] = 52;
razn_w_mem[8557] = 52;
razn_w_mem[8558] = 52;
razn_w_mem[8559] = 52;
razn_w_mem[8560] = 52;
razn_w_mem[8561] = 52;
razn_w_mem[8562] = 52;
razn_w_mem[8563] = 52;
razn_w_mem[8564] = 52;
razn_w_mem[8565] = 52;
razn_w_mem[8566] = 52;
razn_w_mem[8567] = 52;
razn_w_mem[8568] = 52;
razn_w_mem[8569] = 52;
razn_w_mem[8570] = 52;
razn_w_mem[8571] = 52;
razn_w_mem[8572] = 52;
razn_w_mem[8573] = 52;
razn_w_mem[8574] = 52;
razn_w_mem[8575] = 52;
razn_w_mem[8576] = 22;
razn_w_mem[8577] = 22;
razn_w_mem[8578] = 22;
razn_w_mem[8579] = 22;
razn_w_mem[8580] = 22;
razn_w_mem[8581] = 22;
razn_w_mem[8582] = 22;
razn_w_mem[8583] = 22;
razn_w_mem[8584] = 22;
razn_w_mem[8585] = 22;
razn_w_mem[8586] = 22;
razn_w_mem[8587] = 22;
razn_w_mem[8588] = 22;
razn_w_mem[8589] = 22;
razn_w_mem[8590] = 22;
razn_w_mem[8591] = 22;
razn_w_mem[8592] = 22;
razn_w_mem[8593] = 22;
razn_w_mem[8594] = 22;
razn_w_mem[8595] = 22;
razn_w_mem[8596] = 22;
razn_w_mem[8597] = 22;
razn_w_mem[8598] = 22;
razn_w_mem[8599] = 22;
razn_w_mem[8600] = 22;
razn_w_mem[8601] = 22;
razn_w_mem[8602] = 22;
razn_w_mem[8603] = 22;
razn_w_mem[8604] = 22;
razn_w_mem[8605] = 22;
razn_w_mem[8606] = 22;
razn_w_mem[8607] = 22;
razn_w_mem[8608] = 22;
razn_w_mem[8609] = 22;
razn_w_mem[8610] = 22;
razn_w_mem[8611] = 22;
razn_w_mem[8612] = 22;
razn_w_mem[8613] = 22;
razn_w_mem[8614] = 22;
razn_w_mem[8615] = 22;
razn_w_mem[8616] = 22;
razn_w_mem[8617] = 22;
razn_w_mem[8618] = 22;
razn_w_mem[8619] = 22;
razn_w_mem[8620] = 22;
razn_w_mem[8621] = 22;
razn_w_mem[8622] = 22;
razn_w_mem[8623] = 22;
razn_w_mem[8624] = 22;
razn_w_mem[8625] = 22;
razn_w_mem[8626] = 22;
razn_w_mem[8627] = 22;
razn_w_mem[8628] = 22;
razn_w_mem[8629] = 22;
razn_w_mem[8630] = 22;
razn_w_mem[8631] = 22;
razn_w_mem[8632] = 22;
razn_w_mem[8633] = 22;
razn_w_mem[8634] = 22;
razn_w_mem[8635] = 22;
razn_w_mem[8636] = 22;
razn_w_mem[8637] = 22;
razn_w_mem[8638] = 22;
razn_w_mem[8639] = 22;
razn_w_mem[8640] = 22;
razn_w_mem[8641] = 22;
razn_w_mem[8642] = 22;
razn_w_mem[8643] = 22;
razn_w_mem[8644] = 22;
razn_w_mem[8645] = 22;
razn_w_mem[8646] = 22;
razn_w_mem[8647] = 22;
razn_w_mem[8648] = 22;
razn_w_mem[8649] = 22;
razn_w_mem[8650] = 22;
razn_w_mem[8651] = 22;
razn_w_mem[8652] = 22;
razn_w_mem[8653] = 22;
razn_w_mem[8654] = 22;
razn_w_mem[8655] = 22;
razn_w_mem[8656] = 22;
razn_w_mem[8657] = 22;
razn_w_mem[8658] = 22;
razn_w_mem[8659] = 22;
razn_w_mem[8660] = 22;
razn_w_mem[8661] = 22;
razn_w_mem[8662] = 22;
razn_w_mem[8663] = 22;
razn_w_mem[8664] = 22;
razn_w_mem[8665] = 22;
razn_w_mem[8666] = 22;
razn_w_mem[8667] = 22;
razn_w_mem[8668] = 22;
razn_w_mem[8669] = 22;
razn_w_mem[8670] = 22;
razn_w_mem[8671] = 22;
razn_w_mem[8672] = 22;
razn_w_mem[8673] = 22;
razn_w_mem[8674] = 22;
razn_w_mem[8675] = 22;
razn_w_mem[8676] = 22;
razn_w_mem[8677] = 22;
razn_w_mem[8678] = 22;
razn_w_mem[8679] = 22;
razn_w_mem[8680] = 22;
razn_w_mem[8681] = 22;
razn_w_mem[8682] = 22;
razn_w_mem[8683] = 22;
razn_w_mem[8684] = 22;
razn_w_mem[8685] = 22;
razn_w_mem[8686] = 22;
razn_w_mem[8687] = 22;
razn_w_mem[8688] = 22;
razn_w_mem[8689] = 22;
razn_w_mem[8690] = 22;
razn_w_mem[8691] = 22;
razn_w_mem[8692] = 22;
razn_w_mem[8693] = 22;
razn_w_mem[8694] = 22;
razn_w_mem[8695] = 22;
razn_w_mem[8696] = 22;
razn_w_mem[8697] = 22;
razn_w_mem[8698] = 22;
razn_w_mem[8699] = 22;
razn_w_mem[8700] = 22;
razn_w_mem[8701] = 22;
razn_w_mem[8702] = 22;
razn_w_mem[8703] = 22;
razn_w_mem[8704] = 246;
razn_w_mem[8705] = 246;
razn_w_mem[8706] = 246;
razn_w_mem[8707] = 246;
razn_w_mem[8708] = 246;
razn_w_mem[8709] = 246;
razn_w_mem[8710] = 246;
razn_w_mem[8711] = 246;
razn_w_mem[8712] = 246;
razn_w_mem[8713] = 246;
razn_w_mem[8714] = 246;
razn_w_mem[8715] = 246;
razn_w_mem[8716] = 246;
razn_w_mem[8717] = 246;
razn_w_mem[8718] = 246;
razn_w_mem[8719] = 246;
razn_w_mem[8720] = 246;
razn_w_mem[8721] = 246;
razn_w_mem[8722] = 246;
razn_w_mem[8723] = 246;
razn_w_mem[8724] = 246;
razn_w_mem[8725] = 246;
razn_w_mem[8726] = 246;
razn_w_mem[8727] = 246;
razn_w_mem[8728] = 246;
razn_w_mem[8729] = 246;
razn_w_mem[8730] = 246;
razn_w_mem[8731] = 246;
razn_w_mem[8732] = 246;
razn_w_mem[8733] = 246;
razn_w_mem[8734] = 246;
razn_w_mem[8735] = 246;
razn_w_mem[8736] = 246;
razn_w_mem[8737] = 246;
razn_w_mem[8738] = 246;
razn_w_mem[8739] = 246;
razn_w_mem[8740] = 246;
razn_w_mem[8741] = 246;
razn_w_mem[8742] = 246;
razn_w_mem[8743] = 246;
razn_w_mem[8744] = 246;
razn_w_mem[8745] = 246;
razn_w_mem[8746] = 246;
razn_w_mem[8747] = 246;
razn_w_mem[8748] = 246;
razn_w_mem[8749] = 246;
razn_w_mem[8750] = 246;
razn_w_mem[8751] = 246;
razn_w_mem[8752] = 246;
razn_w_mem[8753] = 246;
razn_w_mem[8754] = 246;
razn_w_mem[8755] = 246;
razn_w_mem[8756] = 246;
razn_w_mem[8757] = 246;
razn_w_mem[8758] = 246;
razn_w_mem[8759] = 246;
razn_w_mem[8760] = 246;
razn_w_mem[8761] = 246;
razn_w_mem[8762] = 246;
razn_w_mem[8763] = 246;
razn_w_mem[8764] = 246;
razn_w_mem[8765] = 246;
razn_w_mem[8766] = 246;
razn_w_mem[8767] = 246;
razn_w_mem[8768] = 246;
razn_w_mem[8769] = 246;
razn_w_mem[8770] = 246;
razn_w_mem[8771] = 246;
razn_w_mem[8772] = 246;
razn_w_mem[8773] = 246;
razn_w_mem[8774] = 246;
razn_w_mem[8775] = 246;
razn_w_mem[8776] = 246;
razn_w_mem[8777] = 246;
razn_w_mem[8778] = 246;
razn_w_mem[8779] = 246;
razn_w_mem[8780] = 246;
razn_w_mem[8781] = 246;
razn_w_mem[8782] = 246;
razn_w_mem[8783] = 246;
razn_w_mem[8784] = 246;
razn_w_mem[8785] = 246;
razn_w_mem[8786] = 246;
razn_w_mem[8787] = 246;
razn_w_mem[8788] = 246;
razn_w_mem[8789] = 246;
razn_w_mem[8790] = 246;
razn_w_mem[8791] = 246;
razn_w_mem[8792] = 246;
razn_w_mem[8793] = 246;
razn_w_mem[8794] = 246;
razn_w_mem[8795] = 246;
razn_w_mem[8796] = 246;
razn_w_mem[8797] = 246;
razn_w_mem[8798] = 246;
razn_w_mem[8799] = 246;
razn_w_mem[8800] = 246;
razn_w_mem[8801] = 246;
razn_w_mem[8802] = 246;
razn_w_mem[8803] = 246;
razn_w_mem[8804] = 246;
razn_w_mem[8805] = 246;
razn_w_mem[8806] = 246;
razn_w_mem[8807] = 246;
razn_w_mem[8808] = 246;
razn_w_mem[8809] = 246;
razn_w_mem[8810] = 246;
razn_w_mem[8811] = 246;
razn_w_mem[8812] = 246;
razn_w_mem[8813] = 246;
razn_w_mem[8814] = 246;
razn_w_mem[8815] = 246;
razn_w_mem[8816] = 246;
razn_w_mem[8817] = 246;
razn_w_mem[8818] = 246;
razn_w_mem[8819] = 246;
razn_w_mem[8820] = 246;
razn_w_mem[8821] = 246;
razn_w_mem[8822] = 246;
razn_w_mem[8823] = 246;
razn_w_mem[8824] = 246;
razn_w_mem[8825] = 246;
razn_w_mem[8826] = 246;
razn_w_mem[8827] = 246;
razn_w_mem[8828] = 246;
razn_w_mem[8829] = 246;
razn_w_mem[8830] = 246;
razn_w_mem[8831] = 246;
razn_w_mem[8832] = 216;
razn_w_mem[8833] = 216;
razn_w_mem[8834] = 216;
razn_w_mem[8835] = 216;
razn_w_mem[8836] = 216;
razn_w_mem[8837] = 216;
razn_w_mem[8838] = 216;
razn_w_mem[8839] = 216;
razn_w_mem[8840] = 216;
razn_w_mem[8841] = 216;
razn_w_mem[8842] = 216;
razn_w_mem[8843] = 216;
razn_w_mem[8844] = 216;
razn_w_mem[8845] = 216;
razn_w_mem[8846] = 216;
razn_w_mem[8847] = 216;
razn_w_mem[8848] = 216;
razn_w_mem[8849] = 216;
razn_w_mem[8850] = 216;
razn_w_mem[8851] = 216;
razn_w_mem[8852] = 216;
razn_w_mem[8853] = 216;
razn_w_mem[8854] = 216;
razn_w_mem[8855] = 216;
razn_w_mem[8856] = 216;
razn_w_mem[8857] = 216;
razn_w_mem[8858] = 216;
razn_w_mem[8859] = 216;
razn_w_mem[8860] = 216;
razn_w_mem[8861] = 216;
razn_w_mem[8862] = 216;
razn_w_mem[8863] = 216;
razn_w_mem[8864] = 216;
razn_w_mem[8865] = 216;
razn_w_mem[8866] = 216;
razn_w_mem[8867] = 216;
razn_w_mem[8868] = 216;
razn_w_mem[8869] = 216;
razn_w_mem[8870] = 216;
razn_w_mem[8871] = 216;
razn_w_mem[8872] = 216;
razn_w_mem[8873] = 216;
razn_w_mem[8874] = 216;
razn_w_mem[8875] = 216;
razn_w_mem[8876] = 216;
razn_w_mem[8877] = 216;
razn_w_mem[8878] = 216;
razn_w_mem[8879] = 216;
razn_w_mem[8880] = 216;
razn_w_mem[8881] = 216;
razn_w_mem[8882] = 216;
razn_w_mem[8883] = 216;
razn_w_mem[8884] = 216;
razn_w_mem[8885] = 216;
razn_w_mem[8886] = 216;
razn_w_mem[8887] = 216;
razn_w_mem[8888] = 216;
razn_w_mem[8889] = 216;
razn_w_mem[8890] = 216;
razn_w_mem[8891] = 216;
razn_w_mem[8892] = 216;
razn_w_mem[8893] = 216;
razn_w_mem[8894] = 216;
razn_w_mem[8895] = 216;
razn_w_mem[8896] = 216;
razn_w_mem[8897] = 216;
razn_w_mem[8898] = 216;
razn_w_mem[8899] = 216;
razn_w_mem[8900] = 216;
razn_w_mem[8901] = 216;
razn_w_mem[8902] = 216;
razn_w_mem[8903] = 216;
razn_w_mem[8904] = 216;
razn_w_mem[8905] = 216;
razn_w_mem[8906] = 216;
razn_w_mem[8907] = 216;
razn_w_mem[8908] = 216;
razn_w_mem[8909] = 216;
razn_w_mem[8910] = 216;
razn_w_mem[8911] = 216;
razn_w_mem[8912] = 216;
razn_w_mem[8913] = 216;
razn_w_mem[8914] = 216;
razn_w_mem[8915] = 216;
razn_w_mem[8916] = 216;
razn_w_mem[8917] = 216;
razn_w_mem[8918] = 216;
razn_w_mem[8919] = 216;
razn_w_mem[8920] = 216;
razn_w_mem[8921] = 216;
razn_w_mem[8922] = 216;
razn_w_mem[8923] = 216;
razn_w_mem[8924] = 216;
razn_w_mem[8925] = 216;
razn_w_mem[8926] = 216;
razn_w_mem[8927] = 216;
razn_w_mem[8928] = 216;
razn_w_mem[8929] = 216;
razn_w_mem[8930] = 216;
razn_w_mem[8931] = 216;
razn_w_mem[8932] = 216;
razn_w_mem[8933] = 216;
razn_w_mem[8934] = 216;
razn_w_mem[8935] = 216;
razn_w_mem[8936] = 216;
razn_w_mem[8937] = 216;
razn_w_mem[8938] = 216;
razn_w_mem[8939] = 216;
razn_w_mem[8940] = 216;
razn_w_mem[8941] = 216;
razn_w_mem[8942] = 216;
razn_w_mem[8943] = 216;
razn_w_mem[8944] = 216;
razn_w_mem[8945] = 216;
razn_w_mem[8946] = 216;
razn_w_mem[8947] = 216;
razn_w_mem[8948] = 216;
razn_w_mem[8949] = 216;
razn_w_mem[8950] = 216;
razn_w_mem[8951] = 216;
razn_w_mem[8952] = 216;
razn_w_mem[8953] = 216;
razn_w_mem[8954] = 216;
razn_w_mem[8955] = 216;
razn_w_mem[8956] = 216;
razn_w_mem[8957] = 216;
razn_w_mem[8958] = 216;
razn_w_mem[8959] = 216;
razn_w_mem[8960] = 186;
razn_w_mem[8961] = 186;
razn_w_mem[8962] = 186;
razn_w_mem[8963] = 186;
razn_w_mem[8964] = 186;
razn_w_mem[8965] = 186;
razn_w_mem[8966] = 186;
razn_w_mem[8967] = 186;
razn_w_mem[8968] = 186;
razn_w_mem[8969] = 186;
razn_w_mem[8970] = 186;
razn_w_mem[8971] = 186;
razn_w_mem[8972] = 186;
razn_w_mem[8973] = 186;
razn_w_mem[8974] = 186;
razn_w_mem[8975] = 186;
razn_w_mem[8976] = 186;
razn_w_mem[8977] = 186;
razn_w_mem[8978] = 186;
razn_w_mem[8979] = 186;
razn_w_mem[8980] = 186;
razn_w_mem[8981] = 186;
razn_w_mem[8982] = 186;
razn_w_mem[8983] = 186;
razn_w_mem[8984] = 186;
razn_w_mem[8985] = 186;
razn_w_mem[8986] = 186;
razn_w_mem[8987] = 186;
razn_w_mem[8988] = 186;
razn_w_mem[8989] = 186;
razn_w_mem[8990] = 186;
razn_w_mem[8991] = 186;
razn_w_mem[8992] = 186;
razn_w_mem[8993] = 186;
razn_w_mem[8994] = 186;
razn_w_mem[8995] = 186;
razn_w_mem[8996] = 186;
razn_w_mem[8997] = 186;
razn_w_mem[8998] = 186;
razn_w_mem[8999] = 186;
razn_w_mem[9000] = 186;
razn_w_mem[9001] = 186;
razn_w_mem[9002] = 186;
razn_w_mem[9003] = 186;
razn_w_mem[9004] = 186;
razn_w_mem[9005] = 186;
razn_w_mem[9006] = 186;
razn_w_mem[9007] = 186;
razn_w_mem[9008] = 186;
razn_w_mem[9009] = 186;
razn_w_mem[9010] = 186;
razn_w_mem[9011] = 186;
razn_w_mem[9012] = 186;
razn_w_mem[9013] = 186;
razn_w_mem[9014] = 186;
razn_w_mem[9015] = 186;
razn_w_mem[9016] = 186;
razn_w_mem[9017] = 186;
razn_w_mem[9018] = 186;
razn_w_mem[9019] = 186;
razn_w_mem[9020] = 186;
razn_w_mem[9021] = 186;
razn_w_mem[9022] = 186;
razn_w_mem[9023] = 186;
razn_w_mem[9024] = 186;
razn_w_mem[9025] = 186;
razn_w_mem[9026] = 186;
razn_w_mem[9027] = 186;
razn_w_mem[9028] = 186;
razn_w_mem[9029] = 186;
razn_w_mem[9030] = 186;
razn_w_mem[9031] = 186;
razn_w_mem[9032] = 186;
razn_w_mem[9033] = 186;
razn_w_mem[9034] = 186;
razn_w_mem[9035] = 186;
razn_w_mem[9036] = 186;
razn_w_mem[9037] = 186;
razn_w_mem[9038] = 186;
razn_w_mem[9039] = 186;
razn_w_mem[9040] = 186;
razn_w_mem[9041] = 186;
razn_w_mem[9042] = 186;
razn_w_mem[9043] = 186;
razn_w_mem[9044] = 186;
razn_w_mem[9045] = 186;
razn_w_mem[9046] = 186;
razn_w_mem[9047] = 186;
razn_w_mem[9048] = 186;
razn_w_mem[9049] = 186;
razn_w_mem[9050] = 186;
razn_w_mem[9051] = 186;
razn_w_mem[9052] = 186;
razn_w_mem[9053] = 186;
razn_w_mem[9054] = 186;
razn_w_mem[9055] = 186;
razn_w_mem[9056] = 186;
razn_w_mem[9057] = 186;
razn_w_mem[9058] = 186;
razn_w_mem[9059] = 186;
razn_w_mem[9060] = 186;
razn_w_mem[9061] = 186;
razn_w_mem[9062] = 186;
razn_w_mem[9063] = 186;
razn_w_mem[9064] = 186;
razn_w_mem[9065] = 186;
razn_w_mem[9066] = 186;
razn_w_mem[9067] = 186;
razn_w_mem[9068] = 186;
razn_w_mem[9069] = 186;
razn_w_mem[9070] = 186;
razn_w_mem[9071] = 186;
razn_w_mem[9072] = 186;
razn_w_mem[9073] = 186;
razn_w_mem[9074] = 186;
razn_w_mem[9075] = 186;
razn_w_mem[9076] = 186;
razn_w_mem[9077] = 186;
razn_w_mem[9078] = 186;
razn_w_mem[9079] = 186;
razn_w_mem[9080] = 186;
razn_w_mem[9081] = 186;
razn_w_mem[9082] = 186;
razn_w_mem[9083] = 186;
razn_w_mem[9084] = 186;
razn_w_mem[9085] = 186;
razn_w_mem[9086] = 186;
razn_w_mem[9087] = 186;
razn_w_mem[9088] = 156;
razn_w_mem[9089] = 156;
razn_w_mem[9090] = 156;
razn_w_mem[9091] = 156;
razn_w_mem[9092] = 156;
razn_w_mem[9093] = 156;
razn_w_mem[9094] = 156;
razn_w_mem[9095] = 156;
razn_w_mem[9096] = 156;
razn_w_mem[9097] = 156;
razn_w_mem[9098] = 156;
razn_w_mem[9099] = 156;
razn_w_mem[9100] = 156;
razn_w_mem[9101] = 156;
razn_w_mem[9102] = 156;
razn_w_mem[9103] = 156;
razn_w_mem[9104] = 156;
razn_w_mem[9105] = 156;
razn_w_mem[9106] = 156;
razn_w_mem[9107] = 156;
razn_w_mem[9108] = 156;
razn_w_mem[9109] = 156;
razn_w_mem[9110] = 156;
razn_w_mem[9111] = 156;
razn_w_mem[9112] = 156;
razn_w_mem[9113] = 156;
razn_w_mem[9114] = 156;
razn_w_mem[9115] = 156;
razn_w_mem[9116] = 156;
razn_w_mem[9117] = 156;
razn_w_mem[9118] = 156;
razn_w_mem[9119] = 156;
razn_w_mem[9120] = 156;
razn_w_mem[9121] = 156;
razn_w_mem[9122] = 156;
razn_w_mem[9123] = 156;
razn_w_mem[9124] = 156;
razn_w_mem[9125] = 156;
razn_w_mem[9126] = 156;
razn_w_mem[9127] = 156;
razn_w_mem[9128] = 156;
razn_w_mem[9129] = 156;
razn_w_mem[9130] = 156;
razn_w_mem[9131] = 156;
razn_w_mem[9132] = 156;
razn_w_mem[9133] = 156;
razn_w_mem[9134] = 156;
razn_w_mem[9135] = 156;
razn_w_mem[9136] = 156;
razn_w_mem[9137] = 156;
razn_w_mem[9138] = 156;
razn_w_mem[9139] = 156;
razn_w_mem[9140] = 156;
razn_w_mem[9141] = 156;
razn_w_mem[9142] = 156;
razn_w_mem[9143] = 156;
razn_w_mem[9144] = 156;
razn_w_mem[9145] = 156;
razn_w_mem[9146] = 156;
razn_w_mem[9147] = 156;
razn_w_mem[9148] = 156;
razn_w_mem[9149] = 156;
razn_w_mem[9150] = 156;
razn_w_mem[9151] = 156;
razn_w_mem[9152] = 156;
razn_w_mem[9153] = 156;
razn_w_mem[9154] = 156;
razn_w_mem[9155] = 156;
razn_w_mem[9156] = 156;
razn_w_mem[9157] = 156;
razn_w_mem[9158] = 156;
razn_w_mem[9159] = 156;
razn_w_mem[9160] = 156;
razn_w_mem[9161] = 156;
razn_w_mem[9162] = 156;
razn_w_mem[9163] = 156;
razn_w_mem[9164] = 156;
razn_w_mem[9165] = 156;
razn_w_mem[9166] = 156;
razn_w_mem[9167] = 156;
razn_w_mem[9168] = 156;
razn_w_mem[9169] = 156;
razn_w_mem[9170] = 156;
razn_w_mem[9171] = 156;
razn_w_mem[9172] = 156;
razn_w_mem[9173] = 156;
razn_w_mem[9174] = 156;
razn_w_mem[9175] = 156;
razn_w_mem[9176] = 156;
razn_w_mem[9177] = 156;
razn_w_mem[9178] = 156;
razn_w_mem[9179] = 156;
razn_w_mem[9180] = 156;
razn_w_mem[9181] = 156;
razn_w_mem[9182] = 156;
razn_w_mem[9183] = 156;
razn_w_mem[9184] = 156;
razn_w_mem[9185] = 156;
razn_w_mem[9186] = 156;
razn_w_mem[9187] = 156;
razn_w_mem[9188] = 156;
razn_w_mem[9189] = 156;
razn_w_mem[9190] = 156;
razn_w_mem[9191] = 156;
razn_w_mem[9192] = 156;
razn_w_mem[9193] = 156;
razn_w_mem[9194] = 156;
razn_w_mem[9195] = 156;
razn_w_mem[9196] = 156;
razn_w_mem[9197] = 156;
razn_w_mem[9198] = 156;
razn_w_mem[9199] = 156;
razn_w_mem[9200] = 156;
razn_w_mem[9201] = 156;
razn_w_mem[9202] = 156;
razn_w_mem[9203] = 156;
razn_w_mem[9204] = 156;
razn_w_mem[9205] = 156;
razn_w_mem[9206] = 156;
razn_w_mem[9207] = 156;
razn_w_mem[9208] = 156;
razn_w_mem[9209] = 156;
razn_w_mem[9210] = 156;
razn_w_mem[9211] = 156;
razn_w_mem[9212] = 156;
razn_w_mem[9213] = 156;
razn_w_mem[9214] = 156;
razn_w_mem[9215] = 156;
razn_w_mem[9216] = 126;
razn_w_mem[9217] = 126;
razn_w_mem[9218] = 126;
razn_w_mem[9219] = 126;
razn_w_mem[9220] = 126;
razn_w_mem[9221] = 126;
razn_w_mem[9222] = 126;
razn_w_mem[9223] = 126;
razn_w_mem[9224] = 126;
razn_w_mem[9225] = 126;
razn_w_mem[9226] = 126;
razn_w_mem[9227] = 126;
razn_w_mem[9228] = 126;
razn_w_mem[9229] = 126;
razn_w_mem[9230] = 126;
razn_w_mem[9231] = 126;
razn_w_mem[9232] = 126;
razn_w_mem[9233] = 126;
razn_w_mem[9234] = 126;
razn_w_mem[9235] = 126;
razn_w_mem[9236] = 126;
razn_w_mem[9237] = 126;
razn_w_mem[9238] = 126;
razn_w_mem[9239] = 126;
razn_w_mem[9240] = 126;
razn_w_mem[9241] = 126;
razn_w_mem[9242] = 126;
razn_w_mem[9243] = 126;
razn_w_mem[9244] = 126;
razn_w_mem[9245] = 126;
razn_w_mem[9246] = 126;
razn_w_mem[9247] = 126;
razn_w_mem[9248] = 126;
razn_w_mem[9249] = 126;
razn_w_mem[9250] = 126;
razn_w_mem[9251] = 126;
razn_w_mem[9252] = 126;
razn_w_mem[9253] = 126;
razn_w_mem[9254] = 126;
razn_w_mem[9255] = 126;
razn_w_mem[9256] = 126;
razn_w_mem[9257] = 126;
razn_w_mem[9258] = 126;
razn_w_mem[9259] = 126;
razn_w_mem[9260] = 126;
razn_w_mem[9261] = 126;
razn_w_mem[9262] = 126;
razn_w_mem[9263] = 126;
razn_w_mem[9264] = 126;
razn_w_mem[9265] = 126;
razn_w_mem[9266] = 126;
razn_w_mem[9267] = 126;
razn_w_mem[9268] = 126;
razn_w_mem[9269] = 126;
razn_w_mem[9270] = 126;
razn_w_mem[9271] = 126;
razn_w_mem[9272] = 126;
razn_w_mem[9273] = 126;
razn_w_mem[9274] = 126;
razn_w_mem[9275] = 126;
razn_w_mem[9276] = 126;
razn_w_mem[9277] = 126;
razn_w_mem[9278] = 126;
razn_w_mem[9279] = 126;
razn_w_mem[9280] = 126;
razn_w_mem[9281] = 126;
razn_w_mem[9282] = 126;
razn_w_mem[9283] = 126;
razn_w_mem[9284] = 126;
razn_w_mem[9285] = 126;
razn_w_mem[9286] = 126;
razn_w_mem[9287] = 126;
razn_w_mem[9288] = 126;
razn_w_mem[9289] = 126;
razn_w_mem[9290] = 126;
razn_w_mem[9291] = 126;
razn_w_mem[9292] = 126;
razn_w_mem[9293] = 126;
razn_w_mem[9294] = 126;
razn_w_mem[9295] = 126;
razn_w_mem[9296] = 126;
razn_w_mem[9297] = 126;
razn_w_mem[9298] = 126;
razn_w_mem[9299] = 126;
razn_w_mem[9300] = 126;
razn_w_mem[9301] = 126;
razn_w_mem[9302] = 126;
razn_w_mem[9303] = 126;
razn_w_mem[9304] = 126;
razn_w_mem[9305] = 126;
razn_w_mem[9306] = 126;
razn_w_mem[9307] = 126;
razn_w_mem[9308] = 126;
razn_w_mem[9309] = 126;
razn_w_mem[9310] = 126;
razn_w_mem[9311] = 126;
razn_w_mem[9312] = 126;
razn_w_mem[9313] = 126;
razn_w_mem[9314] = 126;
razn_w_mem[9315] = 126;
razn_w_mem[9316] = 126;
razn_w_mem[9317] = 126;
razn_w_mem[9318] = 126;
razn_w_mem[9319] = 126;
razn_w_mem[9320] = 126;
razn_w_mem[9321] = 126;
razn_w_mem[9322] = 126;
razn_w_mem[9323] = 126;
razn_w_mem[9324] = 126;
razn_w_mem[9325] = 126;
razn_w_mem[9326] = 126;
razn_w_mem[9327] = 126;
razn_w_mem[9328] = 126;
razn_w_mem[9329] = 126;
razn_w_mem[9330] = 126;
razn_w_mem[9331] = 126;
razn_w_mem[9332] = 126;
razn_w_mem[9333] = 126;
razn_w_mem[9334] = 126;
razn_w_mem[9335] = 126;
razn_w_mem[9336] = 126;
razn_w_mem[9337] = 126;
razn_w_mem[9338] = 126;
razn_w_mem[9339] = 126;
razn_w_mem[9340] = 126;
razn_w_mem[9341] = 126;
razn_w_mem[9342] = 126;
razn_w_mem[9343] = 126;
razn_w_mem[9344] = 96;
razn_w_mem[9345] = 96;
razn_w_mem[9346] = 96;
razn_w_mem[9347] = 96;
razn_w_mem[9348] = 96;
razn_w_mem[9349] = 96;
razn_w_mem[9350] = 96;
razn_w_mem[9351] = 96;
razn_w_mem[9352] = 96;
razn_w_mem[9353] = 96;
razn_w_mem[9354] = 96;
razn_w_mem[9355] = 96;
razn_w_mem[9356] = 96;
razn_w_mem[9357] = 96;
razn_w_mem[9358] = 96;
razn_w_mem[9359] = 96;
razn_w_mem[9360] = 96;
razn_w_mem[9361] = 96;
razn_w_mem[9362] = 96;
razn_w_mem[9363] = 96;
razn_w_mem[9364] = 96;
razn_w_mem[9365] = 96;
razn_w_mem[9366] = 96;
razn_w_mem[9367] = 96;
razn_w_mem[9368] = 96;
razn_w_mem[9369] = 96;
razn_w_mem[9370] = 96;
razn_w_mem[9371] = 96;
razn_w_mem[9372] = 96;
razn_w_mem[9373] = 96;
razn_w_mem[9374] = 96;
razn_w_mem[9375] = 96;
razn_w_mem[9376] = 96;
razn_w_mem[9377] = 96;
razn_w_mem[9378] = 96;
razn_w_mem[9379] = 96;
razn_w_mem[9380] = 96;
razn_w_mem[9381] = 96;
razn_w_mem[9382] = 96;
razn_w_mem[9383] = 96;
razn_w_mem[9384] = 96;
razn_w_mem[9385] = 96;
razn_w_mem[9386] = 96;
razn_w_mem[9387] = 96;
razn_w_mem[9388] = 96;
razn_w_mem[9389] = 96;
razn_w_mem[9390] = 96;
razn_w_mem[9391] = 96;
razn_w_mem[9392] = 96;
razn_w_mem[9393] = 96;
razn_w_mem[9394] = 96;
razn_w_mem[9395] = 96;
razn_w_mem[9396] = 96;
razn_w_mem[9397] = 96;
razn_w_mem[9398] = 96;
razn_w_mem[9399] = 96;
razn_w_mem[9400] = 96;
razn_w_mem[9401] = 96;
razn_w_mem[9402] = 96;
razn_w_mem[9403] = 96;
razn_w_mem[9404] = 96;
razn_w_mem[9405] = 96;
razn_w_mem[9406] = 96;
razn_w_mem[9407] = 96;
razn_w_mem[9408] = 96;
razn_w_mem[9409] = 96;
razn_w_mem[9410] = 96;
razn_w_mem[9411] = 96;
razn_w_mem[9412] = 96;
razn_w_mem[9413] = 96;
razn_w_mem[9414] = 96;
razn_w_mem[9415] = 96;
razn_w_mem[9416] = 96;
razn_w_mem[9417] = 96;
razn_w_mem[9418] = 96;
razn_w_mem[9419] = 96;
razn_w_mem[9420] = 96;
razn_w_mem[9421] = 96;
razn_w_mem[9422] = 96;
razn_w_mem[9423] = 96;
razn_w_mem[9424] = 96;
razn_w_mem[9425] = 96;
razn_w_mem[9426] = 96;
razn_w_mem[9427] = 96;
razn_w_mem[9428] = 96;
razn_w_mem[9429] = 96;
razn_w_mem[9430] = 96;
razn_w_mem[9431] = 96;
razn_w_mem[9432] = 96;
razn_w_mem[9433] = 96;
razn_w_mem[9434] = 96;
razn_w_mem[9435] = 96;
razn_w_mem[9436] = 96;
razn_w_mem[9437] = 96;
razn_w_mem[9438] = 96;
razn_w_mem[9439] = 96;
razn_w_mem[9440] = 96;
razn_w_mem[9441] = 96;
razn_w_mem[9442] = 96;
razn_w_mem[9443] = 96;
razn_w_mem[9444] = 96;
razn_w_mem[9445] = 96;
razn_w_mem[9446] = 96;
razn_w_mem[9447] = 96;
razn_w_mem[9448] = 96;
razn_w_mem[9449] = 96;
razn_w_mem[9450] = 96;
razn_w_mem[9451] = 96;
razn_w_mem[9452] = 96;
razn_w_mem[9453] = 96;
razn_w_mem[9454] = 96;
razn_w_mem[9455] = 96;
razn_w_mem[9456] = 96;
razn_w_mem[9457] = 96;
razn_w_mem[9458] = 96;
razn_w_mem[9459] = 96;
razn_w_mem[9460] = 96;
razn_w_mem[9461] = 96;
razn_w_mem[9462] = 96;
razn_w_mem[9463] = 96;
razn_w_mem[9464] = 96;
razn_w_mem[9465] = 96;
razn_w_mem[9466] = 96;
razn_w_mem[9467] = 96;
razn_w_mem[9468] = 96;
razn_w_mem[9469] = 96;
razn_w_mem[9470] = 96;
razn_w_mem[9471] = 96;
razn_w_mem[9472] = 66;
razn_w_mem[9473] = 66;
razn_w_mem[9474] = 66;
razn_w_mem[9475] = 66;
razn_w_mem[9476] = 66;
razn_w_mem[9477] = 66;
razn_w_mem[9478] = 66;
razn_w_mem[9479] = 66;
razn_w_mem[9480] = 66;
razn_w_mem[9481] = 66;
razn_w_mem[9482] = 66;
razn_w_mem[9483] = 66;
razn_w_mem[9484] = 66;
razn_w_mem[9485] = 66;
razn_w_mem[9486] = 66;
razn_w_mem[9487] = 66;
razn_w_mem[9488] = 66;
razn_w_mem[9489] = 66;
razn_w_mem[9490] = 66;
razn_w_mem[9491] = 66;
razn_w_mem[9492] = 66;
razn_w_mem[9493] = 66;
razn_w_mem[9494] = 66;
razn_w_mem[9495] = 66;
razn_w_mem[9496] = 66;
razn_w_mem[9497] = 66;
razn_w_mem[9498] = 66;
razn_w_mem[9499] = 66;
razn_w_mem[9500] = 66;
razn_w_mem[9501] = 66;
razn_w_mem[9502] = 66;
razn_w_mem[9503] = 66;
razn_w_mem[9504] = 66;
razn_w_mem[9505] = 66;
razn_w_mem[9506] = 66;
razn_w_mem[9507] = 66;
razn_w_mem[9508] = 66;
razn_w_mem[9509] = 66;
razn_w_mem[9510] = 66;
razn_w_mem[9511] = 66;
razn_w_mem[9512] = 66;
razn_w_mem[9513] = 66;
razn_w_mem[9514] = 66;
razn_w_mem[9515] = 66;
razn_w_mem[9516] = 66;
razn_w_mem[9517] = 66;
razn_w_mem[9518] = 66;
razn_w_mem[9519] = 66;
razn_w_mem[9520] = 66;
razn_w_mem[9521] = 66;
razn_w_mem[9522] = 66;
razn_w_mem[9523] = 66;
razn_w_mem[9524] = 66;
razn_w_mem[9525] = 66;
razn_w_mem[9526] = 66;
razn_w_mem[9527] = 66;
razn_w_mem[9528] = 66;
razn_w_mem[9529] = 66;
razn_w_mem[9530] = 66;
razn_w_mem[9531] = 66;
razn_w_mem[9532] = 66;
razn_w_mem[9533] = 66;
razn_w_mem[9534] = 66;
razn_w_mem[9535] = 66;
razn_w_mem[9536] = 66;
razn_w_mem[9537] = 66;
razn_w_mem[9538] = 66;
razn_w_mem[9539] = 66;
razn_w_mem[9540] = 66;
razn_w_mem[9541] = 66;
razn_w_mem[9542] = 66;
razn_w_mem[9543] = 66;
razn_w_mem[9544] = 66;
razn_w_mem[9545] = 66;
razn_w_mem[9546] = 66;
razn_w_mem[9547] = 66;
razn_w_mem[9548] = 66;
razn_w_mem[9549] = 66;
razn_w_mem[9550] = 66;
razn_w_mem[9551] = 66;
razn_w_mem[9552] = 66;
razn_w_mem[9553] = 66;
razn_w_mem[9554] = 66;
razn_w_mem[9555] = 66;
razn_w_mem[9556] = 66;
razn_w_mem[9557] = 66;
razn_w_mem[9558] = 66;
razn_w_mem[9559] = 66;
razn_w_mem[9560] = 66;
razn_w_mem[9561] = 66;
razn_w_mem[9562] = 66;
razn_w_mem[9563] = 66;
razn_w_mem[9564] = 66;
razn_w_mem[9565] = 66;
razn_w_mem[9566] = 66;
razn_w_mem[9567] = 66;
razn_w_mem[9568] = 66;
razn_w_mem[9569] = 66;
razn_w_mem[9570] = 66;
razn_w_mem[9571] = 66;
razn_w_mem[9572] = 66;
razn_w_mem[9573] = 66;
razn_w_mem[9574] = 66;
razn_w_mem[9575] = 66;
razn_w_mem[9576] = 66;
razn_w_mem[9577] = 66;
razn_w_mem[9578] = 66;
razn_w_mem[9579] = 66;
razn_w_mem[9580] = 66;
razn_w_mem[9581] = 66;
razn_w_mem[9582] = 66;
razn_w_mem[9583] = 66;
razn_w_mem[9584] = 66;
razn_w_mem[9585] = 66;
razn_w_mem[9586] = 66;
razn_w_mem[9587] = 66;
razn_w_mem[9588] = 66;
razn_w_mem[9589] = 66;
razn_w_mem[9590] = 66;
razn_w_mem[9591] = 66;
razn_w_mem[9592] = 66;
razn_w_mem[9593] = 66;
razn_w_mem[9594] = 66;
razn_w_mem[9595] = 66;
razn_w_mem[9596] = 66;
razn_w_mem[9597] = 66;
razn_w_mem[9598] = 66;
razn_w_mem[9599] = 66;
razn_w_mem[9600] = 36;
razn_w_mem[9601] = 36;
razn_w_mem[9602] = 36;
razn_w_mem[9603] = 36;
razn_w_mem[9604] = 36;
razn_w_mem[9605] = 36;
razn_w_mem[9606] = 36;
razn_w_mem[9607] = 36;
razn_w_mem[9608] = 36;
razn_w_mem[9609] = 36;
razn_w_mem[9610] = 36;
razn_w_mem[9611] = 36;
razn_w_mem[9612] = 36;
razn_w_mem[9613] = 36;
razn_w_mem[9614] = 36;
razn_w_mem[9615] = 36;
razn_w_mem[9616] = 36;
razn_w_mem[9617] = 36;
razn_w_mem[9618] = 36;
razn_w_mem[9619] = 36;
razn_w_mem[9620] = 36;
razn_w_mem[9621] = 36;
razn_w_mem[9622] = 36;
razn_w_mem[9623] = 36;
razn_w_mem[9624] = 36;
razn_w_mem[9625] = 36;
razn_w_mem[9626] = 36;
razn_w_mem[9627] = 36;
razn_w_mem[9628] = 36;
razn_w_mem[9629] = 36;
razn_w_mem[9630] = 36;
razn_w_mem[9631] = 36;
razn_w_mem[9632] = 36;
razn_w_mem[9633] = 36;
razn_w_mem[9634] = 36;
razn_w_mem[9635] = 36;
razn_w_mem[9636] = 36;
razn_w_mem[9637] = 36;
razn_w_mem[9638] = 36;
razn_w_mem[9639] = 36;
razn_w_mem[9640] = 36;
razn_w_mem[9641] = 36;
razn_w_mem[9642] = 36;
razn_w_mem[9643] = 36;
razn_w_mem[9644] = 36;
razn_w_mem[9645] = 36;
razn_w_mem[9646] = 36;
razn_w_mem[9647] = 36;
razn_w_mem[9648] = 36;
razn_w_mem[9649] = 36;
razn_w_mem[9650] = 36;
razn_w_mem[9651] = 36;
razn_w_mem[9652] = 36;
razn_w_mem[9653] = 36;
razn_w_mem[9654] = 36;
razn_w_mem[9655] = 36;
razn_w_mem[9656] = 36;
razn_w_mem[9657] = 36;
razn_w_mem[9658] = 36;
razn_w_mem[9659] = 36;
razn_w_mem[9660] = 36;
razn_w_mem[9661] = 36;
razn_w_mem[9662] = 36;
razn_w_mem[9663] = 36;
razn_w_mem[9664] = 36;
razn_w_mem[9665] = 36;
razn_w_mem[9666] = 36;
razn_w_mem[9667] = 36;
razn_w_mem[9668] = 36;
razn_w_mem[9669] = 36;
razn_w_mem[9670] = 36;
razn_w_mem[9671] = 36;
razn_w_mem[9672] = 36;
razn_w_mem[9673] = 36;
razn_w_mem[9674] = 36;
razn_w_mem[9675] = 36;
razn_w_mem[9676] = 36;
razn_w_mem[9677] = 36;
razn_w_mem[9678] = 36;
razn_w_mem[9679] = 36;
razn_w_mem[9680] = 36;
razn_w_mem[9681] = 36;
razn_w_mem[9682] = 36;
razn_w_mem[9683] = 36;
razn_w_mem[9684] = 36;
razn_w_mem[9685] = 36;
razn_w_mem[9686] = 36;
razn_w_mem[9687] = 36;
razn_w_mem[9688] = 36;
razn_w_mem[9689] = 36;
razn_w_mem[9690] = 36;
razn_w_mem[9691] = 36;
razn_w_mem[9692] = 36;
razn_w_mem[9693] = 36;
razn_w_mem[9694] = 36;
razn_w_mem[9695] = 36;
razn_w_mem[9696] = 36;
razn_w_mem[9697] = 36;
razn_w_mem[9698] = 36;
razn_w_mem[9699] = 36;
razn_w_mem[9700] = 36;
razn_w_mem[9701] = 36;
razn_w_mem[9702] = 36;
razn_w_mem[9703] = 36;
razn_w_mem[9704] = 36;
razn_w_mem[9705] = 36;
razn_w_mem[9706] = 36;
razn_w_mem[9707] = 36;
razn_w_mem[9708] = 36;
razn_w_mem[9709] = 36;
razn_w_mem[9710] = 36;
razn_w_mem[9711] = 36;
razn_w_mem[9712] = 36;
razn_w_mem[9713] = 36;
razn_w_mem[9714] = 36;
razn_w_mem[9715] = 36;
razn_w_mem[9716] = 36;
razn_w_mem[9717] = 36;
razn_w_mem[9718] = 36;
razn_w_mem[9719] = 36;
razn_w_mem[9720] = 36;
razn_w_mem[9721] = 36;
razn_w_mem[9722] = 36;
razn_w_mem[9723] = 36;
razn_w_mem[9724] = 36;
razn_w_mem[9725] = 36;
razn_w_mem[9726] = 36;
razn_w_mem[9727] = 36;
razn_w_mem[9728] = 6;
razn_w_mem[9729] = 6;
razn_w_mem[9730] = 6;
razn_w_mem[9731] = 6;
razn_w_mem[9732] = 6;
razn_w_mem[9733] = 6;
razn_w_mem[9734] = 6;
razn_w_mem[9735] = 6;
razn_w_mem[9736] = 6;
razn_w_mem[9737] = 6;
razn_w_mem[9738] = 6;
razn_w_mem[9739] = 6;
razn_w_mem[9740] = 6;
razn_w_mem[9741] = 6;
razn_w_mem[9742] = 6;
razn_w_mem[9743] = 6;
razn_w_mem[9744] = 6;
razn_w_mem[9745] = 6;
razn_w_mem[9746] = 6;
razn_w_mem[9747] = 6;
razn_w_mem[9748] = 6;
razn_w_mem[9749] = 6;
razn_w_mem[9750] = 6;
razn_w_mem[9751] = 6;
razn_w_mem[9752] = 6;
razn_w_mem[9753] = 6;
razn_w_mem[9754] = 6;
razn_w_mem[9755] = 6;
razn_w_mem[9756] = 6;
razn_w_mem[9757] = 6;
razn_w_mem[9758] = 6;
razn_w_mem[9759] = 6;
razn_w_mem[9760] = 6;
razn_w_mem[9761] = 6;
razn_w_mem[9762] = 6;
razn_w_mem[9763] = 6;
razn_w_mem[9764] = 6;
razn_w_mem[9765] = 6;
razn_w_mem[9766] = 6;
razn_w_mem[9767] = 6;
razn_w_mem[9768] = 6;
razn_w_mem[9769] = 6;
razn_w_mem[9770] = 6;
razn_w_mem[9771] = 6;
razn_w_mem[9772] = 6;
razn_w_mem[9773] = 6;
razn_w_mem[9774] = 6;
razn_w_mem[9775] = 6;
razn_w_mem[9776] = 6;
razn_w_mem[9777] = 6;
razn_w_mem[9778] = 6;
razn_w_mem[9779] = 6;
razn_w_mem[9780] = 6;
razn_w_mem[9781] = 6;
razn_w_mem[9782] = 6;
razn_w_mem[9783] = 6;
razn_w_mem[9784] = 6;
razn_w_mem[9785] = 6;
razn_w_mem[9786] = 6;
razn_w_mem[9787] = 6;
razn_w_mem[9788] = 6;
razn_w_mem[9789] = 6;
razn_w_mem[9790] = 6;
razn_w_mem[9791] = 6;
razn_w_mem[9792] = 6;
razn_w_mem[9793] = 6;
razn_w_mem[9794] = 6;
razn_w_mem[9795] = 6;
razn_w_mem[9796] = 6;
razn_w_mem[9797] = 6;
razn_w_mem[9798] = 6;
razn_w_mem[9799] = 6;
razn_w_mem[9800] = 6;
razn_w_mem[9801] = 6;
razn_w_mem[9802] = 6;
razn_w_mem[9803] = 6;
razn_w_mem[9804] = 6;
razn_w_mem[9805] = 6;
razn_w_mem[9806] = 6;
razn_w_mem[9807] = 6;
razn_w_mem[9808] = 6;
razn_w_mem[9809] = 6;
razn_w_mem[9810] = 6;
razn_w_mem[9811] = 6;
razn_w_mem[9812] = 6;
razn_w_mem[9813] = 6;
razn_w_mem[9814] = 6;
razn_w_mem[9815] = 6;
razn_w_mem[9816] = 6;
razn_w_mem[9817] = 6;
razn_w_mem[9818] = 6;
razn_w_mem[9819] = 6;
razn_w_mem[9820] = 6;
razn_w_mem[9821] = 6;
razn_w_mem[9822] = 6;
razn_w_mem[9823] = 6;
razn_w_mem[9824] = 6;
razn_w_mem[9825] = 6;
razn_w_mem[9826] = 6;
razn_w_mem[9827] = 6;
razn_w_mem[9828] = 6;
razn_w_mem[9829] = 6;
razn_w_mem[9830] = 6;
razn_w_mem[9831] = 6;
razn_w_mem[9832] = 6;
razn_w_mem[9833] = 6;
razn_w_mem[9834] = 6;
razn_w_mem[9835] = 6;
razn_w_mem[9836] = 6;
razn_w_mem[9837] = 6;
razn_w_mem[9838] = 6;
razn_w_mem[9839] = 6;
razn_w_mem[9840] = 6;
razn_w_mem[9841] = 6;
razn_w_mem[9842] = 6;
razn_w_mem[9843] = 6;
razn_w_mem[9844] = 6;
razn_w_mem[9845] = 6;
razn_w_mem[9846] = 6;
razn_w_mem[9847] = 6;
razn_w_mem[9848] = 6;
razn_w_mem[9849] = 6;
razn_w_mem[9850] = 6;
razn_w_mem[9851] = 6;
razn_w_mem[9852] = 6;
razn_w_mem[9853] = 6;
razn_w_mem[9854] = 6;
razn_w_mem[9855] = 6;
razn_w_mem[9856] = 230;
razn_w_mem[9857] = 230;
razn_w_mem[9858] = 230;
razn_w_mem[9859] = 230;
razn_w_mem[9860] = 230;
razn_w_mem[9861] = 230;
razn_w_mem[9862] = 230;
razn_w_mem[9863] = 230;
razn_w_mem[9864] = 230;
razn_w_mem[9865] = 230;
razn_w_mem[9866] = 230;
razn_w_mem[9867] = 230;
razn_w_mem[9868] = 230;
razn_w_mem[9869] = 230;
razn_w_mem[9870] = 230;
razn_w_mem[9871] = 230;
razn_w_mem[9872] = 230;
razn_w_mem[9873] = 230;
razn_w_mem[9874] = 230;
razn_w_mem[9875] = 230;
razn_w_mem[9876] = 230;
razn_w_mem[9877] = 230;
razn_w_mem[9878] = 230;
razn_w_mem[9879] = 230;
razn_w_mem[9880] = 230;
razn_w_mem[9881] = 230;
razn_w_mem[9882] = 230;
razn_w_mem[9883] = 230;
razn_w_mem[9884] = 230;
razn_w_mem[9885] = 230;
razn_w_mem[9886] = 230;
razn_w_mem[9887] = 230;
razn_w_mem[9888] = 230;
razn_w_mem[9889] = 230;
razn_w_mem[9890] = 230;
razn_w_mem[9891] = 230;
razn_w_mem[9892] = 230;
razn_w_mem[9893] = 230;
razn_w_mem[9894] = 230;
razn_w_mem[9895] = 230;
razn_w_mem[9896] = 230;
razn_w_mem[9897] = 230;
razn_w_mem[9898] = 230;
razn_w_mem[9899] = 230;
razn_w_mem[9900] = 230;
razn_w_mem[9901] = 230;
razn_w_mem[9902] = 230;
razn_w_mem[9903] = 230;
razn_w_mem[9904] = 230;
razn_w_mem[9905] = 230;
razn_w_mem[9906] = 230;
razn_w_mem[9907] = 230;
razn_w_mem[9908] = 230;
razn_w_mem[9909] = 230;
razn_w_mem[9910] = 230;
razn_w_mem[9911] = 230;
razn_w_mem[9912] = 230;
razn_w_mem[9913] = 230;
razn_w_mem[9914] = 230;
razn_w_mem[9915] = 230;
razn_w_mem[9916] = 230;
razn_w_mem[9917] = 230;
razn_w_mem[9918] = 230;
razn_w_mem[9919] = 230;
razn_w_mem[9920] = 230;
razn_w_mem[9921] = 230;
razn_w_mem[9922] = 230;
razn_w_mem[9923] = 230;
razn_w_mem[9924] = 230;
razn_w_mem[9925] = 230;
razn_w_mem[9926] = 230;
razn_w_mem[9927] = 230;
razn_w_mem[9928] = 230;
razn_w_mem[9929] = 230;
razn_w_mem[9930] = 230;
razn_w_mem[9931] = 230;
razn_w_mem[9932] = 230;
razn_w_mem[9933] = 230;
razn_w_mem[9934] = 230;
razn_w_mem[9935] = 230;
razn_w_mem[9936] = 230;
razn_w_mem[9937] = 230;
razn_w_mem[9938] = 230;
razn_w_mem[9939] = 230;
razn_w_mem[9940] = 230;
razn_w_mem[9941] = 230;
razn_w_mem[9942] = 230;
razn_w_mem[9943] = 230;
razn_w_mem[9944] = 230;
razn_w_mem[9945] = 230;
razn_w_mem[9946] = 230;
razn_w_mem[9947] = 230;
razn_w_mem[9948] = 230;
razn_w_mem[9949] = 230;
razn_w_mem[9950] = 230;
razn_w_mem[9951] = 230;
razn_w_mem[9952] = 230;
razn_w_mem[9953] = 230;
razn_w_mem[9954] = 230;
razn_w_mem[9955] = 230;
razn_w_mem[9956] = 230;
razn_w_mem[9957] = 230;
razn_w_mem[9958] = 230;
razn_w_mem[9959] = 230;
razn_w_mem[9960] = 230;
razn_w_mem[9961] = 230;
razn_w_mem[9962] = 230;
razn_w_mem[9963] = 230;
razn_w_mem[9964] = 230;
razn_w_mem[9965] = 230;
razn_w_mem[9966] = 230;
razn_w_mem[9967] = 230;
razn_w_mem[9968] = 230;
razn_w_mem[9969] = 230;
razn_w_mem[9970] = 230;
razn_w_mem[9971] = 230;
razn_w_mem[9972] = 230;
razn_w_mem[9973] = 230;
razn_w_mem[9974] = 230;
razn_w_mem[9975] = 230;
razn_w_mem[9976] = 230;
razn_w_mem[9977] = 230;
razn_w_mem[9978] = 230;
razn_w_mem[9979] = 230;
razn_w_mem[9980] = 230;
razn_w_mem[9981] = 230;
razn_w_mem[9982] = 230;
razn_w_mem[9983] = 230;
razn_w_mem[9984] = 200;
razn_w_mem[9985] = 200;
razn_w_mem[9986] = 200;
razn_w_mem[9987] = 200;
razn_w_mem[9988] = 200;
razn_w_mem[9989] = 200;
razn_w_mem[9990] = 200;
razn_w_mem[9991] = 200;
razn_w_mem[9992] = 200;
razn_w_mem[9993] = 200;
razn_w_mem[9994] = 200;
razn_w_mem[9995] = 200;
razn_w_mem[9996] = 200;
razn_w_mem[9997] = 200;
razn_w_mem[9998] = 200;
razn_w_mem[9999] = 200;
razn_w_mem[10000] = 200;
razn_w_mem[10001] = 200;
razn_w_mem[10002] = 200;
razn_w_mem[10003] = 200;
razn_w_mem[10004] = 200;
razn_w_mem[10005] = 200;
razn_w_mem[10006] = 200;
razn_w_mem[10007] = 200;
razn_w_mem[10008] = 200;
razn_w_mem[10009] = 200;
razn_w_mem[10010] = 200;
razn_w_mem[10011] = 200;
razn_w_mem[10012] = 200;
razn_w_mem[10013] = 200;
razn_w_mem[10014] = 200;
razn_w_mem[10015] = 200;
razn_w_mem[10016] = 200;
razn_w_mem[10017] = 200;
razn_w_mem[10018] = 200;
razn_w_mem[10019] = 200;
razn_w_mem[10020] = 200;
razn_w_mem[10021] = 200;
razn_w_mem[10022] = 200;
razn_w_mem[10023] = 200;
razn_w_mem[10024] = 200;
razn_w_mem[10025] = 200;
razn_w_mem[10026] = 200;
razn_w_mem[10027] = 200;
razn_w_mem[10028] = 200;
razn_w_mem[10029] = 200;
razn_w_mem[10030] = 200;
razn_w_mem[10031] = 200;
razn_w_mem[10032] = 200;
razn_w_mem[10033] = 200;
razn_w_mem[10034] = 200;
razn_w_mem[10035] = 200;
razn_w_mem[10036] = 200;
razn_w_mem[10037] = 200;
razn_w_mem[10038] = 200;
razn_w_mem[10039] = 200;
razn_w_mem[10040] = 200;
razn_w_mem[10041] = 200;
razn_w_mem[10042] = 200;
razn_w_mem[10043] = 200;
razn_w_mem[10044] = 200;
razn_w_mem[10045] = 200;
razn_w_mem[10046] = 200;
razn_w_mem[10047] = 200;
razn_w_mem[10048] = 200;
razn_w_mem[10049] = 200;
razn_w_mem[10050] = 200;
razn_w_mem[10051] = 200;
razn_w_mem[10052] = 200;
razn_w_mem[10053] = 200;
razn_w_mem[10054] = 200;
razn_w_mem[10055] = 200;
razn_w_mem[10056] = 200;
razn_w_mem[10057] = 200;
razn_w_mem[10058] = 200;
razn_w_mem[10059] = 200;
razn_w_mem[10060] = 200;
razn_w_mem[10061] = 200;
razn_w_mem[10062] = 200;
razn_w_mem[10063] = 200;
razn_w_mem[10064] = 200;
razn_w_mem[10065] = 200;
razn_w_mem[10066] = 200;
razn_w_mem[10067] = 200;
razn_w_mem[10068] = 200;
razn_w_mem[10069] = 200;
razn_w_mem[10070] = 200;
razn_w_mem[10071] = 200;
razn_w_mem[10072] = 200;
razn_w_mem[10073] = 200;
razn_w_mem[10074] = 200;
razn_w_mem[10075] = 200;
razn_w_mem[10076] = 200;
razn_w_mem[10077] = 200;
razn_w_mem[10078] = 200;
razn_w_mem[10079] = 200;
razn_w_mem[10080] = 200;
razn_w_mem[10081] = 200;
razn_w_mem[10082] = 200;
razn_w_mem[10083] = 200;
razn_w_mem[10084] = 200;
razn_w_mem[10085] = 200;
razn_w_mem[10086] = 200;
razn_w_mem[10087] = 200;
razn_w_mem[10088] = 200;
razn_w_mem[10089] = 200;
razn_w_mem[10090] = 200;
razn_w_mem[10091] = 200;
razn_w_mem[10092] = 200;
razn_w_mem[10093] = 200;
razn_w_mem[10094] = 200;
razn_w_mem[10095] = 200;
razn_w_mem[10096] = 200;
razn_w_mem[10097] = 200;
razn_w_mem[10098] = 200;
razn_w_mem[10099] = 200;
razn_w_mem[10100] = 200;
razn_w_mem[10101] = 200;
razn_w_mem[10102] = 200;
razn_w_mem[10103] = 200;
razn_w_mem[10104] = 200;
razn_w_mem[10105] = 200;
razn_w_mem[10106] = 200;
razn_w_mem[10107] = 200;
razn_w_mem[10108] = 200;
razn_w_mem[10109] = 200;
razn_w_mem[10110] = 200;
razn_w_mem[10111] = 200;
razn_w_mem[10112] = 170;
razn_w_mem[10113] = 170;
razn_w_mem[10114] = 170;
razn_w_mem[10115] = 170;
razn_w_mem[10116] = 170;
razn_w_mem[10117] = 170;
razn_w_mem[10118] = 170;
razn_w_mem[10119] = 170;
razn_w_mem[10120] = 170;
razn_w_mem[10121] = 170;
razn_w_mem[10122] = 170;
razn_w_mem[10123] = 170;
razn_w_mem[10124] = 170;
razn_w_mem[10125] = 170;
razn_w_mem[10126] = 170;
razn_w_mem[10127] = 170;
razn_w_mem[10128] = 170;
razn_w_mem[10129] = 170;
razn_w_mem[10130] = 170;
razn_w_mem[10131] = 170;
razn_w_mem[10132] = 170;
razn_w_mem[10133] = 170;
razn_w_mem[10134] = 170;
razn_w_mem[10135] = 170;
razn_w_mem[10136] = 170;
razn_w_mem[10137] = 170;
razn_w_mem[10138] = 170;
razn_w_mem[10139] = 170;
razn_w_mem[10140] = 170;
razn_w_mem[10141] = 170;
razn_w_mem[10142] = 170;
razn_w_mem[10143] = 170;
razn_w_mem[10144] = 170;
razn_w_mem[10145] = 170;
razn_w_mem[10146] = 170;
razn_w_mem[10147] = 170;
razn_w_mem[10148] = 170;
razn_w_mem[10149] = 170;
razn_w_mem[10150] = 170;
razn_w_mem[10151] = 170;
razn_w_mem[10152] = 170;
razn_w_mem[10153] = 170;
razn_w_mem[10154] = 170;
razn_w_mem[10155] = 170;
razn_w_mem[10156] = 170;
razn_w_mem[10157] = 170;
razn_w_mem[10158] = 170;
razn_w_mem[10159] = 170;
razn_w_mem[10160] = 170;
razn_w_mem[10161] = 170;
razn_w_mem[10162] = 170;
razn_w_mem[10163] = 170;
razn_w_mem[10164] = 170;
razn_w_mem[10165] = 170;
razn_w_mem[10166] = 170;
razn_w_mem[10167] = 170;
razn_w_mem[10168] = 170;
razn_w_mem[10169] = 170;
razn_w_mem[10170] = 170;
razn_w_mem[10171] = 170;
razn_w_mem[10172] = 170;
razn_w_mem[10173] = 170;
razn_w_mem[10174] = 170;
razn_w_mem[10175] = 170;
razn_w_mem[10176] = 170;
razn_w_mem[10177] = 170;
razn_w_mem[10178] = 170;
razn_w_mem[10179] = 170;
razn_w_mem[10180] = 170;
razn_w_mem[10181] = 170;
razn_w_mem[10182] = 170;
razn_w_mem[10183] = 170;
razn_w_mem[10184] = 170;
razn_w_mem[10185] = 170;
razn_w_mem[10186] = 170;
razn_w_mem[10187] = 170;
razn_w_mem[10188] = 170;
razn_w_mem[10189] = 170;
razn_w_mem[10190] = 170;
razn_w_mem[10191] = 170;
razn_w_mem[10192] = 170;
razn_w_mem[10193] = 170;
razn_w_mem[10194] = 170;
razn_w_mem[10195] = 170;
razn_w_mem[10196] = 170;
razn_w_mem[10197] = 170;
razn_w_mem[10198] = 170;
razn_w_mem[10199] = 170;
razn_w_mem[10200] = 170;
razn_w_mem[10201] = 170;
razn_w_mem[10202] = 170;
razn_w_mem[10203] = 170;
razn_w_mem[10204] = 170;
razn_w_mem[10205] = 170;
razn_w_mem[10206] = 170;
razn_w_mem[10207] = 170;
razn_w_mem[10208] = 170;
razn_w_mem[10209] = 170;
razn_w_mem[10210] = 170;
razn_w_mem[10211] = 170;
razn_w_mem[10212] = 170;
razn_w_mem[10213] = 170;
razn_w_mem[10214] = 170;
razn_w_mem[10215] = 170;
razn_w_mem[10216] = 170;
razn_w_mem[10217] = 170;
razn_w_mem[10218] = 170;
razn_w_mem[10219] = 170;
razn_w_mem[10220] = 170;
razn_w_mem[10221] = 170;
razn_w_mem[10222] = 170;
razn_w_mem[10223] = 170;
razn_w_mem[10224] = 170;
razn_w_mem[10225] = 170;
razn_w_mem[10226] = 170;
razn_w_mem[10227] = 170;
razn_w_mem[10228] = 170;
razn_w_mem[10229] = 170;
razn_w_mem[10230] = 170;
razn_w_mem[10231] = 170;
razn_w_mem[10232] = 170;
razn_w_mem[10233] = 170;
razn_w_mem[10234] = 170;
razn_w_mem[10235] = 170;
razn_w_mem[10236] = 170;
razn_w_mem[10237] = 170;
razn_w_mem[10238] = 170;
razn_w_mem[10239] = 170;
razn_w_mem[10240] = 140;
razn_w_mem[10241] = 140;
razn_w_mem[10242] = 140;
razn_w_mem[10243] = 140;
razn_w_mem[10244] = 140;
razn_w_mem[10245] = 140;
razn_w_mem[10246] = 140;
razn_w_mem[10247] = 140;
razn_w_mem[10248] = 140;
razn_w_mem[10249] = 140;
razn_w_mem[10250] = 140;
razn_w_mem[10251] = 140;
razn_w_mem[10252] = 140;
razn_w_mem[10253] = 140;
razn_w_mem[10254] = 140;
razn_w_mem[10255] = 140;
razn_w_mem[10256] = 140;
razn_w_mem[10257] = 140;
razn_w_mem[10258] = 140;
razn_w_mem[10259] = 140;
razn_w_mem[10260] = 140;
razn_w_mem[10261] = 140;
razn_w_mem[10262] = 140;
razn_w_mem[10263] = 140;
razn_w_mem[10264] = 140;
razn_w_mem[10265] = 140;
razn_w_mem[10266] = 140;
razn_w_mem[10267] = 140;
razn_w_mem[10268] = 140;
razn_w_mem[10269] = 140;
razn_w_mem[10270] = 140;
razn_w_mem[10271] = 140;
razn_w_mem[10272] = 140;
razn_w_mem[10273] = 140;
razn_w_mem[10274] = 140;
razn_w_mem[10275] = 140;
razn_w_mem[10276] = 140;
razn_w_mem[10277] = 140;
razn_w_mem[10278] = 140;
razn_w_mem[10279] = 140;
razn_w_mem[10280] = 140;
razn_w_mem[10281] = 140;
razn_w_mem[10282] = 140;
razn_w_mem[10283] = 140;
razn_w_mem[10284] = 140;
razn_w_mem[10285] = 140;
razn_w_mem[10286] = 140;
razn_w_mem[10287] = 140;
razn_w_mem[10288] = 140;
razn_w_mem[10289] = 140;
razn_w_mem[10290] = 140;
razn_w_mem[10291] = 140;
razn_w_mem[10292] = 140;
razn_w_mem[10293] = 140;
razn_w_mem[10294] = 140;
razn_w_mem[10295] = 140;
razn_w_mem[10296] = 140;
razn_w_mem[10297] = 140;
razn_w_mem[10298] = 140;
razn_w_mem[10299] = 140;
razn_w_mem[10300] = 140;
razn_w_mem[10301] = 140;
razn_w_mem[10302] = 140;
razn_w_mem[10303] = 140;
razn_w_mem[10304] = 140;
razn_w_mem[10305] = 140;
razn_w_mem[10306] = 140;
razn_w_mem[10307] = 140;
razn_w_mem[10308] = 140;
razn_w_mem[10309] = 140;
razn_w_mem[10310] = 140;
razn_w_mem[10311] = 140;
razn_w_mem[10312] = 140;
razn_w_mem[10313] = 140;
razn_w_mem[10314] = 140;
razn_w_mem[10315] = 140;
razn_w_mem[10316] = 140;
razn_w_mem[10317] = 140;
razn_w_mem[10318] = 140;
razn_w_mem[10319] = 140;
razn_w_mem[10320] = 140;
razn_w_mem[10321] = 140;
razn_w_mem[10322] = 140;
razn_w_mem[10323] = 140;
razn_w_mem[10324] = 140;
razn_w_mem[10325] = 140;
razn_w_mem[10326] = 140;
razn_w_mem[10327] = 140;
razn_w_mem[10328] = 140;
razn_w_mem[10329] = 140;
razn_w_mem[10330] = 140;
razn_w_mem[10331] = 140;
razn_w_mem[10332] = 140;
razn_w_mem[10333] = 140;
razn_w_mem[10334] = 140;
razn_w_mem[10335] = 140;
razn_w_mem[10336] = 140;
razn_w_mem[10337] = 140;
razn_w_mem[10338] = 140;
razn_w_mem[10339] = 140;
razn_w_mem[10340] = 140;
razn_w_mem[10341] = 140;
razn_w_mem[10342] = 140;
razn_w_mem[10343] = 140;
razn_w_mem[10344] = 140;
razn_w_mem[10345] = 140;
razn_w_mem[10346] = 140;
razn_w_mem[10347] = 140;
razn_w_mem[10348] = 140;
razn_w_mem[10349] = 140;
razn_w_mem[10350] = 140;
razn_w_mem[10351] = 140;
razn_w_mem[10352] = 140;
razn_w_mem[10353] = 140;
razn_w_mem[10354] = 140;
razn_w_mem[10355] = 140;
razn_w_mem[10356] = 140;
razn_w_mem[10357] = 140;
razn_w_mem[10358] = 140;
razn_w_mem[10359] = 140;
razn_w_mem[10360] = 140;
razn_w_mem[10361] = 140;
razn_w_mem[10362] = 140;
razn_w_mem[10363] = 140;
razn_w_mem[10364] = 140;
razn_w_mem[10365] = 140;
razn_w_mem[10366] = 140;
razn_w_mem[10367] = 140;
razn_w_mem[10368] = 110;
razn_w_mem[10369] = 110;
razn_w_mem[10370] = 110;
razn_w_mem[10371] = 110;
razn_w_mem[10372] = 110;
razn_w_mem[10373] = 110;
razn_w_mem[10374] = 110;
razn_w_mem[10375] = 110;
razn_w_mem[10376] = 110;
razn_w_mem[10377] = 110;
razn_w_mem[10378] = 110;
razn_w_mem[10379] = 110;
razn_w_mem[10380] = 110;
razn_w_mem[10381] = 110;
razn_w_mem[10382] = 110;
razn_w_mem[10383] = 110;
razn_w_mem[10384] = 110;
razn_w_mem[10385] = 110;
razn_w_mem[10386] = 110;
razn_w_mem[10387] = 110;
razn_w_mem[10388] = 110;
razn_w_mem[10389] = 110;
razn_w_mem[10390] = 110;
razn_w_mem[10391] = 110;
razn_w_mem[10392] = 110;
razn_w_mem[10393] = 110;
razn_w_mem[10394] = 110;
razn_w_mem[10395] = 110;
razn_w_mem[10396] = 110;
razn_w_mem[10397] = 110;
razn_w_mem[10398] = 110;
razn_w_mem[10399] = 110;
razn_w_mem[10400] = 110;
razn_w_mem[10401] = 110;
razn_w_mem[10402] = 110;
razn_w_mem[10403] = 110;
razn_w_mem[10404] = 110;
razn_w_mem[10405] = 110;
razn_w_mem[10406] = 110;
razn_w_mem[10407] = 110;
razn_w_mem[10408] = 110;
razn_w_mem[10409] = 110;
razn_w_mem[10410] = 110;
razn_w_mem[10411] = 110;
razn_w_mem[10412] = 110;
razn_w_mem[10413] = 110;
razn_w_mem[10414] = 110;
razn_w_mem[10415] = 110;
razn_w_mem[10416] = 110;
razn_w_mem[10417] = 110;
razn_w_mem[10418] = 110;
razn_w_mem[10419] = 110;
razn_w_mem[10420] = 110;
razn_w_mem[10421] = 110;
razn_w_mem[10422] = 110;
razn_w_mem[10423] = 110;
razn_w_mem[10424] = 110;
razn_w_mem[10425] = 110;
razn_w_mem[10426] = 110;
razn_w_mem[10427] = 110;
razn_w_mem[10428] = 110;
razn_w_mem[10429] = 110;
razn_w_mem[10430] = 110;
razn_w_mem[10431] = 110;
razn_w_mem[10432] = 110;
razn_w_mem[10433] = 110;
razn_w_mem[10434] = 110;
razn_w_mem[10435] = 110;
razn_w_mem[10436] = 110;
razn_w_mem[10437] = 110;
razn_w_mem[10438] = 110;
razn_w_mem[10439] = 110;
razn_w_mem[10440] = 110;
razn_w_mem[10441] = 110;
razn_w_mem[10442] = 110;
razn_w_mem[10443] = 110;
razn_w_mem[10444] = 110;
razn_w_mem[10445] = 110;
razn_w_mem[10446] = 110;
razn_w_mem[10447] = 110;
razn_w_mem[10448] = 110;
razn_w_mem[10449] = 110;
razn_w_mem[10450] = 110;
razn_w_mem[10451] = 110;
razn_w_mem[10452] = 110;
razn_w_mem[10453] = 110;
razn_w_mem[10454] = 110;
razn_w_mem[10455] = 110;
razn_w_mem[10456] = 110;
razn_w_mem[10457] = 110;
razn_w_mem[10458] = 110;
razn_w_mem[10459] = 110;
razn_w_mem[10460] = 110;
razn_w_mem[10461] = 110;
razn_w_mem[10462] = 110;
razn_w_mem[10463] = 110;
razn_w_mem[10464] = 110;
razn_w_mem[10465] = 110;
razn_w_mem[10466] = 110;
razn_w_mem[10467] = 110;
razn_w_mem[10468] = 110;
razn_w_mem[10469] = 110;
razn_w_mem[10470] = 110;
razn_w_mem[10471] = 110;
razn_w_mem[10472] = 110;
razn_w_mem[10473] = 110;
razn_w_mem[10474] = 110;
razn_w_mem[10475] = 110;
razn_w_mem[10476] = 110;
razn_w_mem[10477] = 110;
razn_w_mem[10478] = 110;
razn_w_mem[10479] = 110;
razn_w_mem[10480] = 110;
razn_w_mem[10481] = 110;
razn_w_mem[10482] = 110;
razn_w_mem[10483] = 110;
razn_w_mem[10484] = 110;
razn_w_mem[10485] = 110;
razn_w_mem[10486] = 110;
razn_w_mem[10487] = 110;
razn_w_mem[10488] = 110;
razn_w_mem[10489] = 110;
razn_w_mem[10490] = 110;
razn_w_mem[10491] = 110;
razn_w_mem[10492] = 110;
razn_w_mem[10493] = 110;
razn_w_mem[10494] = 110;
razn_w_mem[10495] = 110;
razn_w_mem[10496] = 80;
razn_w_mem[10497] = 80;
razn_w_mem[10498] = 80;
razn_w_mem[10499] = 80;
razn_w_mem[10500] = 80;
razn_w_mem[10501] = 80;
razn_w_mem[10502] = 80;
razn_w_mem[10503] = 80;
razn_w_mem[10504] = 80;
razn_w_mem[10505] = 80;
razn_w_mem[10506] = 80;
razn_w_mem[10507] = 80;
razn_w_mem[10508] = 80;
razn_w_mem[10509] = 80;
razn_w_mem[10510] = 80;
razn_w_mem[10511] = 80;
razn_w_mem[10512] = 80;
razn_w_mem[10513] = 80;
razn_w_mem[10514] = 80;
razn_w_mem[10515] = 80;
razn_w_mem[10516] = 80;
razn_w_mem[10517] = 80;
razn_w_mem[10518] = 80;
razn_w_mem[10519] = 80;
razn_w_mem[10520] = 80;
razn_w_mem[10521] = 80;
razn_w_mem[10522] = 80;
razn_w_mem[10523] = 80;
razn_w_mem[10524] = 80;
razn_w_mem[10525] = 80;
razn_w_mem[10526] = 80;
razn_w_mem[10527] = 80;
razn_w_mem[10528] = 80;
razn_w_mem[10529] = 80;
razn_w_mem[10530] = 80;
razn_w_mem[10531] = 80;
razn_w_mem[10532] = 80;
razn_w_mem[10533] = 80;
razn_w_mem[10534] = 80;
razn_w_mem[10535] = 80;
razn_w_mem[10536] = 80;
razn_w_mem[10537] = 80;
razn_w_mem[10538] = 80;
razn_w_mem[10539] = 80;
razn_w_mem[10540] = 80;
razn_w_mem[10541] = 80;
razn_w_mem[10542] = 80;
razn_w_mem[10543] = 80;
razn_w_mem[10544] = 80;
razn_w_mem[10545] = 80;
razn_w_mem[10546] = 80;
razn_w_mem[10547] = 80;
razn_w_mem[10548] = 80;
razn_w_mem[10549] = 80;
razn_w_mem[10550] = 80;
razn_w_mem[10551] = 80;
razn_w_mem[10552] = 80;
razn_w_mem[10553] = 80;
razn_w_mem[10554] = 80;
razn_w_mem[10555] = 80;
razn_w_mem[10556] = 80;
razn_w_mem[10557] = 80;
razn_w_mem[10558] = 80;
razn_w_mem[10559] = 80;
razn_w_mem[10560] = 80;
razn_w_mem[10561] = 80;
razn_w_mem[10562] = 80;
razn_w_mem[10563] = 80;
razn_w_mem[10564] = 80;
razn_w_mem[10565] = 80;
razn_w_mem[10566] = 80;
razn_w_mem[10567] = 80;
razn_w_mem[10568] = 80;
razn_w_mem[10569] = 80;
razn_w_mem[10570] = 80;
razn_w_mem[10571] = 80;
razn_w_mem[10572] = 80;
razn_w_mem[10573] = 80;
razn_w_mem[10574] = 80;
razn_w_mem[10575] = 80;
razn_w_mem[10576] = 80;
razn_w_mem[10577] = 80;
razn_w_mem[10578] = 80;
razn_w_mem[10579] = 80;
razn_w_mem[10580] = 80;
razn_w_mem[10581] = 80;
razn_w_mem[10582] = 80;
razn_w_mem[10583] = 80;
razn_w_mem[10584] = 80;
razn_w_mem[10585] = 80;
razn_w_mem[10586] = 80;
razn_w_mem[10587] = 80;
razn_w_mem[10588] = 80;
razn_w_mem[10589] = 80;
razn_w_mem[10590] = 80;
razn_w_mem[10591] = 80;
razn_w_mem[10592] = 80;
razn_w_mem[10593] = 80;
razn_w_mem[10594] = 80;
razn_w_mem[10595] = 80;
razn_w_mem[10596] = 80;
razn_w_mem[10597] = 80;
razn_w_mem[10598] = 80;
razn_w_mem[10599] = 80;
razn_w_mem[10600] = 80;
razn_w_mem[10601] = 80;
razn_w_mem[10602] = 80;
razn_w_mem[10603] = 80;
razn_w_mem[10604] = 80;
razn_w_mem[10605] = 80;
razn_w_mem[10606] = 80;
razn_w_mem[10607] = 80;
razn_w_mem[10608] = 80;
razn_w_mem[10609] = 80;
razn_w_mem[10610] = 80;
razn_w_mem[10611] = 80;
razn_w_mem[10612] = 80;
razn_w_mem[10613] = 80;
razn_w_mem[10614] = 80;
razn_w_mem[10615] = 80;
razn_w_mem[10616] = 80;
razn_w_mem[10617] = 80;
razn_w_mem[10618] = 80;
razn_w_mem[10619] = 80;
razn_w_mem[10620] = 80;
razn_w_mem[10621] = 80;
razn_w_mem[10622] = 80;
razn_w_mem[10623] = 80;
razn_w_mem[10624] = 50;
razn_w_mem[10625] = 50;
razn_w_mem[10626] = 50;
razn_w_mem[10627] = 50;
razn_w_mem[10628] = 50;
razn_w_mem[10629] = 50;
razn_w_mem[10630] = 50;
razn_w_mem[10631] = 50;
razn_w_mem[10632] = 50;
razn_w_mem[10633] = 50;
razn_w_mem[10634] = 50;
razn_w_mem[10635] = 50;
razn_w_mem[10636] = 50;
razn_w_mem[10637] = 50;
razn_w_mem[10638] = 50;
razn_w_mem[10639] = 50;
razn_w_mem[10640] = 50;
razn_w_mem[10641] = 50;
razn_w_mem[10642] = 50;
razn_w_mem[10643] = 50;
razn_w_mem[10644] = 50;
razn_w_mem[10645] = 50;
razn_w_mem[10646] = 50;
razn_w_mem[10647] = 50;
razn_w_mem[10648] = 50;
razn_w_mem[10649] = 50;
razn_w_mem[10650] = 50;
razn_w_mem[10651] = 50;
razn_w_mem[10652] = 50;
razn_w_mem[10653] = 50;
razn_w_mem[10654] = 50;
razn_w_mem[10655] = 50;
razn_w_mem[10656] = 50;
razn_w_mem[10657] = 50;
razn_w_mem[10658] = 50;
razn_w_mem[10659] = 50;
razn_w_mem[10660] = 50;
razn_w_mem[10661] = 50;
razn_w_mem[10662] = 50;
razn_w_mem[10663] = 50;
razn_w_mem[10664] = 50;
razn_w_mem[10665] = 50;
razn_w_mem[10666] = 50;
razn_w_mem[10667] = 50;
razn_w_mem[10668] = 50;
razn_w_mem[10669] = 50;
razn_w_mem[10670] = 50;
razn_w_mem[10671] = 50;
razn_w_mem[10672] = 50;
razn_w_mem[10673] = 50;
razn_w_mem[10674] = 50;
razn_w_mem[10675] = 50;
razn_w_mem[10676] = 50;
razn_w_mem[10677] = 50;
razn_w_mem[10678] = 50;
razn_w_mem[10679] = 50;
razn_w_mem[10680] = 50;
razn_w_mem[10681] = 50;
razn_w_mem[10682] = 50;
razn_w_mem[10683] = 50;
razn_w_mem[10684] = 50;
razn_w_mem[10685] = 50;
razn_w_mem[10686] = 50;
razn_w_mem[10687] = 50;
razn_w_mem[10688] = 50;
razn_w_mem[10689] = 50;
razn_w_mem[10690] = 50;
razn_w_mem[10691] = 50;
razn_w_mem[10692] = 50;
razn_w_mem[10693] = 50;
razn_w_mem[10694] = 50;
razn_w_mem[10695] = 50;
razn_w_mem[10696] = 50;
razn_w_mem[10697] = 50;
razn_w_mem[10698] = 50;
razn_w_mem[10699] = 50;
razn_w_mem[10700] = 50;
razn_w_mem[10701] = 50;
razn_w_mem[10702] = 50;
razn_w_mem[10703] = 50;
razn_w_mem[10704] = 50;
razn_w_mem[10705] = 50;
razn_w_mem[10706] = 50;
razn_w_mem[10707] = 50;
razn_w_mem[10708] = 50;
razn_w_mem[10709] = 50;
razn_w_mem[10710] = 50;
razn_w_mem[10711] = 50;
razn_w_mem[10712] = 50;
razn_w_mem[10713] = 50;
razn_w_mem[10714] = 50;
razn_w_mem[10715] = 50;
razn_w_mem[10716] = 50;
razn_w_mem[10717] = 50;
razn_w_mem[10718] = 50;
razn_w_mem[10719] = 50;
razn_w_mem[10720] = 50;
razn_w_mem[10721] = 50;
razn_w_mem[10722] = 50;
razn_w_mem[10723] = 50;
razn_w_mem[10724] = 50;
razn_w_mem[10725] = 50;
razn_w_mem[10726] = 50;
razn_w_mem[10727] = 50;
razn_w_mem[10728] = 50;
razn_w_mem[10729] = 50;
razn_w_mem[10730] = 50;
razn_w_mem[10731] = 50;
razn_w_mem[10732] = 50;
razn_w_mem[10733] = 50;
razn_w_mem[10734] = 50;
razn_w_mem[10735] = 50;
razn_w_mem[10736] = 50;
razn_w_mem[10737] = 50;
razn_w_mem[10738] = 50;
razn_w_mem[10739] = 50;
razn_w_mem[10740] = 50;
razn_w_mem[10741] = 50;
razn_w_mem[10742] = 50;
razn_w_mem[10743] = 50;
razn_w_mem[10744] = 50;
razn_w_mem[10745] = 50;
razn_w_mem[10746] = 50;
razn_w_mem[10747] = 50;
razn_w_mem[10748] = 50;
razn_w_mem[10749] = 50;
razn_w_mem[10750] = 50;
razn_w_mem[10751] = 50;
razn_w_mem[10752] = 20;
razn_w_mem[10753] = 20;
razn_w_mem[10754] = 20;
razn_w_mem[10755] = 20;
razn_w_mem[10756] = 20;
razn_w_mem[10757] = 20;
razn_w_mem[10758] = 20;
razn_w_mem[10759] = 20;
razn_w_mem[10760] = 20;
razn_w_mem[10761] = 20;
razn_w_mem[10762] = 20;
razn_w_mem[10763] = 20;
razn_w_mem[10764] = 20;
razn_w_mem[10765] = 20;
razn_w_mem[10766] = 20;
razn_w_mem[10767] = 20;
razn_w_mem[10768] = 20;
razn_w_mem[10769] = 20;
razn_w_mem[10770] = 20;
razn_w_mem[10771] = 20;
razn_w_mem[10772] = 20;
razn_w_mem[10773] = 20;
razn_w_mem[10774] = 20;
razn_w_mem[10775] = 20;
razn_w_mem[10776] = 20;
razn_w_mem[10777] = 20;
razn_w_mem[10778] = 20;
razn_w_mem[10779] = 20;
razn_w_mem[10780] = 20;
razn_w_mem[10781] = 20;
razn_w_mem[10782] = 20;
razn_w_mem[10783] = 20;
razn_w_mem[10784] = 20;
razn_w_mem[10785] = 20;
razn_w_mem[10786] = 20;
razn_w_mem[10787] = 20;
razn_w_mem[10788] = 20;
razn_w_mem[10789] = 20;
razn_w_mem[10790] = 20;
razn_w_mem[10791] = 20;
razn_w_mem[10792] = 20;
razn_w_mem[10793] = 20;
razn_w_mem[10794] = 20;
razn_w_mem[10795] = 20;
razn_w_mem[10796] = 20;
razn_w_mem[10797] = 20;
razn_w_mem[10798] = 20;
razn_w_mem[10799] = 20;
razn_w_mem[10800] = 20;
razn_w_mem[10801] = 20;
razn_w_mem[10802] = 20;
razn_w_mem[10803] = 20;
razn_w_mem[10804] = 20;
razn_w_mem[10805] = 20;
razn_w_mem[10806] = 20;
razn_w_mem[10807] = 20;
razn_w_mem[10808] = 20;
razn_w_mem[10809] = 20;
razn_w_mem[10810] = 20;
razn_w_mem[10811] = 20;
razn_w_mem[10812] = 20;
razn_w_mem[10813] = 20;
razn_w_mem[10814] = 20;
razn_w_mem[10815] = 20;
razn_w_mem[10816] = 20;
razn_w_mem[10817] = 20;
razn_w_mem[10818] = 20;
razn_w_mem[10819] = 20;
razn_w_mem[10820] = 20;
razn_w_mem[10821] = 20;
razn_w_mem[10822] = 20;
razn_w_mem[10823] = 20;
razn_w_mem[10824] = 20;
razn_w_mem[10825] = 20;
razn_w_mem[10826] = 20;
razn_w_mem[10827] = 20;
razn_w_mem[10828] = 20;
razn_w_mem[10829] = 20;
razn_w_mem[10830] = 20;
razn_w_mem[10831] = 20;
razn_w_mem[10832] = 20;
razn_w_mem[10833] = 20;
razn_w_mem[10834] = 20;
razn_w_mem[10835] = 20;
razn_w_mem[10836] = 20;
razn_w_mem[10837] = 20;
razn_w_mem[10838] = 20;
razn_w_mem[10839] = 20;
razn_w_mem[10840] = 20;
razn_w_mem[10841] = 20;
razn_w_mem[10842] = 20;
razn_w_mem[10843] = 20;
razn_w_mem[10844] = 20;
razn_w_mem[10845] = 20;
razn_w_mem[10846] = 20;
razn_w_mem[10847] = 20;
razn_w_mem[10848] = 20;
razn_w_mem[10849] = 20;
razn_w_mem[10850] = 20;
razn_w_mem[10851] = 20;
razn_w_mem[10852] = 20;
razn_w_mem[10853] = 20;
razn_w_mem[10854] = 20;
razn_w_mem[10855] = 20;
razn_w_mem[10856] = 20;
razn_w_mem[10857] = 20;
razn_w_mem[10858] = 20;
razn_w_mem[10859] = 20;
razn_w_mem[10860] = 20;
razn_w_mem[10861] = 20;
razn_w_mem[10862] = 20;
razn_w_mem[10863] = 20;
razn_w_mem[10864] = 20;
razn_w_mem[10865] = 20;
razn_w_mem[10866] = 20;
razn_w_mem[10867] = 20;
razn_w_mem[10868] = 20;
razn_w_mem[10869] = 20;
razn_w_mem[10870] = 20;
razn_w_mem[10871] = 20;
razn_w_mem[10872] = 20;
razn_w_mem[10873] = 20;
razn_w_mem[10874] = 20;
razn_w_mem[10875] = 20;
razn_w_mem[10876] = 20;
razn_w_mem[10877] = 20;
razn_w_mem[10878] = 20;
razn_w_mem[10879] = 20;
razn_w_mem[10880] = 244;
razn_w_mem[10881] = 244;
razn_w_mem[10882] = 244;
razn_w_mem[10883] = 244;
razn_w_mem[10884] = 244;
razn_w_mem[10885] = 244;
razn_w_mem[10886] = 244;
razn_w_mem[10887] = 244;
razn_w_mem[10888] = 244;
razn_w_mem[10889] = 244;
razn_w_mem[10890] = 244;
razn_w_mem[10891] = 244;
razn_w_mem[10892] = 244;
razn_w_mem[10893] = 244;
razn_w_mem[10894] = 244;
razn_w_mem[10895] = 244;
razn_w_mem[10896] = 244;
razn_w_mem[10897] = 244;
razn_w_mem[10898] = 244;
razn_w_mem[10899] = 244;
razn_w_mem[10900] = 244;
razn_w_mem[10901] = 244;
razn_w_mem[10902] = 244;
razn_w_mem[10903] = 244;
razn_w_mem[10904] = 244;
razn_w_mem[10905] = 244;
razn_w_mem[10906] = 244;
razn_w_mem[10907] = 244;
razn_w_mem[10908] = 244;
razn_w_mem[10909] = 244;
razn_w_mem[10910] = 244;
razn_w_mem[10911] = 244;
razn_w_mem[10912] = 244;
razn_w_mem[10913] = 244;
razn_w_mem[10914] = 244;
razn_w_mem[10915] = 244;
razn_w_mem[10916] = 244;
razn_w_mem[10917] = 244;
razn_w_mem[10918] = 244;
razn_w_mem[10919] = 244;
razn_w_mem[10920] = 244;
razn_w_mem[10921] = 244;
razn_w_mem[10922] = 244;
razn_w_mem[10923] = 244;
razn_w_mem[10924] = 244;
razn_w_mem[10925] = 244;
razn_w_mem[10926] = 244;
razn_w_mem[10927] = 244;
razn_w_mem[10928] = 244;
razn_w_mem[10929] = 244;
razn_w_mem[10930] = 244;
razn_w_mem[10931] = 244;
razn_w_mem[10932] = 244;
razn_w_mem[10933] = 244;
razn_w_mem[10934] = 244;
razn_w_mem[10935] = 244;
razn_w_mem[10936] = 244;
razn_w_mem[10937] = 244;
razn_w_mem[10938] = 244;
razn_w_mem[10939] = 244;
razn_w_mem[10940] = 244;
razn_w_mem[10941] = 244;
razn_w_mem[10942] = 244;
razn_w_mem[10943] = 244;
razn_w_mem[10944] = 244;
razn_w_mem[10945] = 244;
razn_w_mem[10946] = 244;
razn_w_mem[10947] = 244;
razn_w_mem[10948] = 244;
razn_w_mem[10949] = 244;
razn_w_mem[10950] = 244;
razn_w_mem[10951] = 244;
razn_w_mem[10952] = 244;
razn_w_mem[10953] = 244;
razn_w_mem[10954] = 244;
razn_w_mem[10955] = 244;
razn_w_mem[10956] = 244;
razn_w_mem[10957] = 244;
razn_w_mem[10958] = 244;
razn_w_mem[10959] = 244;
razn_w_mem[10960] = 244;
razn_w_mem[10961] = 244;
razn_w_mem[10962] = 244;
razn_w_mem[10963] = 244;
razn_w_mem[10964] = 244;
razn_w_mem[10965] = 244;
razn_w_mem[10966] = 244;
razn_w_mem[10967] = 244;
razn_w_mem[10968] = 244;
razn_w_mem[10969] = 244;
razn_w_mem[10970] = 244;
razn_w_mem[10971] = 244;
razn_w_mem[10972] = 244;
razn_w_mem[10973] = 244;
razn_w_mem[10974] = 244;
razn_w_mem[10975] = 244;
razn_w_mem[10976] = 244;
razn_w_mem[10977] = 244;
razn_w_mem[10978] = 244;
razn_w_mem[10979] = 244;
razn_w_mem[10980] = 244;
razn_w_mem[10981] = 244;
razn_w_mem[10982] = 244;
razn_w_mem[10983] = 244;
razn_w_mem[10984] = 244;
razn_w_mem[10985] = 244;
razn_w_mem[10986] = 244;
razn_w_mem[10987] = 244;
razn_w_mem[10988] = 244;
razn_w_mem[10989] = 244;
razn_w_mem[10990] = 244;
razn_w_mem[10991] = 244;
razn_w_mem[10992] = 244;
razn_w_mem[10993] = 244;
razn_w_mem[10994] = 244;
razn_w_mem[10995] = 244;
razn_w_mem[10996] = 244;
razn_w_mem[10997] = 244;
razn_w_mem[10998] = 244;
razn_w_mem[10999] = 244;
razn_w_mem[11000] = 244;
razn_w_mem[11001] = 244;
razn_w_mem[11002] = 244;
razn_w_mem[11003] = 244;
razn_w_mem[11004] = 244;
razn_w_mem[11005] = 244;
razn_w_mem[11006] = 244;
razn_w_mem[11007] = 244;
razn_w_mem[11008] = 214;
razn_w_mem[11009] = 214;
razn_w_mem[11010] = 214;
razn_w_mem[11011] = 214;
razn_w_mem[11012] = 214;
razn_w_mem[11013] = 214;
razn_w_mem[11014] = 214;
razn_w_mem[11015] = 214;
razn_w_mem[11016] = 214;
razn_w_mem[11017] = 214;
razn_w_mem[11018] = 214;
razn_w_mem[11019] = 214;
razn_w_mem[11020] = 214;
razn_w_mem[11021] = 214;
razn_w_mem[11022] = 214;
razn_w_mem[11023] = 214;
razn_w_mem[11024] = 214;
razn_w_mem[11025] = 214;
razn_w_mem[11026] = 214;
razn_w_mem[11027] = 214;
razn_w_mem[11028] = 214;
razn_w_mem[11029] = 214;
razn_w_mem[11030] = 214;
razn_w_mem[11031] = 214;
razn_w_mem[11032] = 214;
razn_w_mem[11033] = 214;
razn_w_mem[11034] = 214;
razn_w_mem[11035] = 214;
razn_w_mem[11036] = 214;
razn_w_mem[11037] = 214;
razn_w_mem[11038] = 214;
razn_w_mem[11039] = 214;
razn_w_mem[11040] = 214;
razn_w_mem[11041] = 214;
razn_w_mem[11042] = 214;
razn_w_mem[11043] = 214;
razn_w_mem[11044] = 214;
razn_w_mem[11045] = 214;
razn_w_mem[11046] = 214;
razn_w_mem[11047] = 214;
razn_w_mem[11048] = 214;
razn_w_mem[11049] = 214;
razn_w_mem[11050] = 214;
razn_w_mem[11051] = 214;
razn_w_mem[11052] = 214;
razn_w_mem[11053] = 214;
razn_w_mem[11054] = 214;
razn_w_mem[11055] = 214;
razn_w_mem[11056] = 214;
razn_w_mem[11057] = 214;
razn_w_mem[11058] = 214;
razn_w_mem[11059] = 214;
razn_w_mem[11060] = 214;
razn_w_mem[11061] = 214;
razn_w_mem[11062] = 214;
razn_w_mem[11063] = 214;
razn_w_mem[11064] = 214;
razn_w_mem[11065] = 214;
razn_w_mem[11066] = 214;
razn_w_mem[11067] = 214;
razn_w_mem[11068] = 214;
razn_w_mem[11069] = 214;
razn_w_mem[11070] = 214;
razn_w_mem[11071] = 214;
razn_w_mem[11072] = 214;
razn_w_mem[11073] = 214;
razn_w_mem[11074] = 214;
razn_w_mem[11075] = 214;
razn_w_mem[11076] = 214;
razn_w_mem[11077] = 214;
razn_w_mem[11078] = 214;
razn_w_mem[11079] = 214;
razn_w_mem[11080] = 214;
razn_w_mem[11081] = 214;
razn_w_mem[11082] = 214;
razn_w_mem[11083] = 214;
razn_w_mem[11084] = 214;
razn_w_mem[11085] = 214;
razn_w_mem[11086] = 214;
razn_w_mem[11087] = 214;
razn_w_mem[11088] = 214;
razn_w_mem[11089] = 214;
razn_w_mem[11090] = 214;
razn_w_mem[11091] = 214;
razn_w_mem[11092] = 214;
razn_w_mem[11093] = 214;
razn_w_mem[11094] = 214;
razn_w_mem[11095] = 214;
razn_w_mem[11096] = 214;
razn_w_mem[11097] = 214;
razn_w_mem[11098] = 214;
razn_w_mem[11099] = 214;
razn_w_mem[11100] = 214;
razn_w_mem[11101] = 214;
razn_w_mem[11102] = 214;
razn_w_mem[11103] = 214;
razn_w_mem[11104] = 214;
razn_w_mem[11105] = 214;
razn_w_mem[11106] = 214;
razn_w_mem[11107] = 214;
razn_w_mem[11108] = 214;
razn_w_mem[11109] = 214;
razn_w_mem[11110] = 214;
razn_w_mem[11111] = 214;
razn_w_mem[11112] = 214;
razn_w_mem[11113] = 214;
razn_w_mem[11114] = 214;
razn_w_mem[11115] = 214;
razn_w_mem[11116] = 214;
razn_w_mem[11117] = 214;
razn_w_mem[11118] = 214;
razn_w_mem[11119] = 214;
razn_w_mem[11120] = 214;
razn_w_mem[11121] = 214;
razn_w_mem[11122] = 214;
razn_w_mem[11123] = 214;
razn_w_mem[11124] = 214;
razn_w_mem[11125] = 214;
razn_w_mem[11126] = 214;
razn_w_mem[11127] = 214;
razn_w_mem[11128] = 214;
razn_w_mem[11129] = 214;
razn_w_mem[11130] = 214;
razn_w_mem[11131] = 214;
razn_w_mem[11132] = 214;
razn_w_mem[11133] = 214;
razn_w_mem[11134] = 214;
razn_w_mem[11135] = 214;
razn_w_mem[11136] = 184;
razn_w_mem[11137] = 184;
razn_w_mem[11138] = 184;
razn_w_mem[11139] = 184;
razn_w_mem[11140] = 184;
razn_w_mem[11141] = 184;
razn_w_mem[11142] = 184;
razn_w_mem[11143] = 184;
razn_w_mem[11144] = 184;
razn_w_mem[11145] = 184;
razn_w_mem[11146] = 184;
razn_w_mem[11147] = 184;
razn_w_mem[11148] = 184;
razn_w_mem[11149] = 184;
razn_w_mem[11150] = 184;
razn_w_mem[11151] = 184;
razn_w_mem[11152] = 184;
razn_w_mem[11153] = 184;
razn_w_mem[11154] = 184;
razn_w_mem[11155] = 184;
razn_w_mem[11156] = 184;
razn_w_mem[11157] = 184;
razn_w_mem[11158] = 184;
razn_w_mem[11159] = 184;
razn_w_mem[11160] = 184;
razn_w_mem[11161] = 184;
razn_w_mem[11162] = 184;
razn_w_mem[11163] = 184;
razn_w_mem[11164] = 184;
razn_w_mem[11165] = 184;
razn_w_mem[11166] = 184;
razn_w_mem[11167] = 184;
razn_w_mem[11168] = 184;
razn_w_mem[11169] = 184;
razn_w_mem[11170] = 184;
razn_w_mem[11171] = 184;
razn_w_mem[11172] = 184;
razn_w_mem[11173] = 184;
razn_w_mem[11174] = 184;
razn_w_mem[11175] = 184;
razn_w_mem[11176] = 184;
razn_w_mem[11177] = 184;
razn_w_mem[11178] = 184;
razn_w_mem[11179] = 184;
razn_w_mem[11180] = 184;
razn_w_mem[11181] = 184;
razn_w_mem[11182] = 184;
razn_w_mem[11183] = 184;
razn_w_mem[11184] = 184;
razn_w_mem[11185] = 184;
razn_w_mem[11186] = 184;
razn_w_mem[11187] = 184;
razn_w_mem[11188] = 184;
razn_w_mem[11189] = 184;
razn_w_mem[11190] = 184;
razn_w_mem[11191] = 184;
razn_w_mem[11192] = 184;
razn_w_mem[11193] = 184;
razn_w_mem[11194] = 184;
razn_w_mem[11195] = 184;
razn_w_mem[11196] = 184;
razn_w_mem[11197] = 184;
razn_w_mem[11198] = 184;
razn_w_mem[11199] = 184;
razn_w_mem[11200] = 184;
razn_w_mem[11201] = 184;
razn_w_mem[11202] = 184;
razn_w_mem[11203] = 184;
razn_w_mem[11204] = 184;
razn_w_mem[11205] = 184;
razn_w_mem[11206] = 184;
razn_w_mem[11207] = 184;
razn_w_mem[11208] = 184;
razn_w_mem[11209] = 184;
razn_w_mem[11210] = 184;
razn_w_mem[11211] = 184;
razn_w_mem[11212] = 184;
razn_w_mem[11213] = 184;
razn_w_mem[11214] = 184;
razn_w_mem[11215] = 184;
razn_w_mem[11216] = 184;
razn_w_mem[11217] = 184;
razn_w_mem[11218] = 184;
razn_w_mem[11219] = 184;
razn_w_mem[11220] = 184;
razn_w_mem[11221] = 184;
razn_w_mem[11222] = 184;
razn_w_mem[11223] = 184;
razn_w_mem[11224] = 184;
razn_w_mem[11225] = 184;
razn_w_mem[11226] = 184;
razn_w_mem[11227] = 184;
razn_w_mem[11228] = 184;
razn_w_mem[11229] = 184;
razn_w_mem[11230] = 184;
razn_w_mem[11231] = 184;
razn_w_mem[11232] = 184;
razn_w_mem[11233] = 184;
razn_w_mem[11234] = 184;
razn_w_mem[11235] = 184;
razn_w_mem[11236] = 184;
razn_w_mem[11237] = 184;
razn_w_mem[11238] = 184;
razn_w_mem[11239] = 184;
razn_w_mem[11240] = 184;
razn_w_mem[11241] = 184;
razn_w_mem[11242] = 184;
razn_w_mem[11243] = 184;
razn_w_mem[11244] = 184;
razn_w_mem[11245] = 184;
razn_w_mem[11246] = 184;
razn_w_mem[11247] = 184;
razn_w_mem[11248] = 184;
razn_w_mem[11249] = 184;
razn_w_mem[11250] = 184;
razn_w_mem[11251] = 184;
razn_w_mem[11252] = 184;
razn_w_mem[11253] = 184;
razn_w_mem[11254] = 184;
razn_w_mem[11255] = 184;
razn_w_mem[11256] = 184;
razn_w_mem[11257] = 184;
razn_w_mem[11258] = 184;
razn_w_mem[11259] = 184;
razn_w_mem[11260] = 184;
razn_w_mem[11261] = 184;
razn_w_mem[11262] = 184;
razn_w_mem[11263] = 184;
razn_w_mem[11264] = 154;
razn_w_mem[11265] = 154;
razn_w_mem[11266] = 154;
razn_w_mem[11267] = 154;
razn_w_mem[11268] = 154;
razn_w_mem[11269] = 154;
razn_w_mem[11270] = 154;
razn_w_mem[11271] = 154;
razn_w_mem[11272] = 154;
razn_w_mem[11273] = 154;
razn_w_mem[11274] = 154;
razn_w_mem[11275] = 154;
razn_w_mem[11276] = 154;
razn_w_mem[11277] = 154;
razn_w_mem[11278] = 154;
razn_w_mem[11279] = 154;
razn_w_mem[11280] = 154;
razn_w_mem[11281] = 154;
razn_w_mem[11282] = 154;
razn_w_mem[11283] = 154;
razn_w_mem[11284] = 154;
razn_w_mem[11285] = 154;
razn_w_mem[11286] = 154;
razn_w_mem[11287] = 154;
razn_w_mem[11288] = 154;
razn_w_mem[11289] = 154;
razn_w_mem[11290] = 154;
razn_w_mem[11291] = 154;
razn_w_mem[11292] = 154;
razn_w_mem[11293] = 154;
razn_w_mem[11294] = 154;
razn_w_mem[11295] = 154;
razn_w_mem[11296] = 154;
razn_w_mem[11297] = 154;
razn_w_mem[11298] = 154;
razn_w_mem[11299] = 154;
razn_w_mem[11300] = 154;
razn_w_mem[11301] = 154;
razn_w_mem[11302] = 154;
razn_w_mem[11303] = 154;
razn_w_mem[11304] = 154;
razn_w_mem[11305] = 154;
razn_w_mem[11306] = 154;
razn_w_mem[11307] = 154;
razn_w_mem[11308] = 154;
razn_w_mem[11309] = 154;
razn_w_mem[11310] = 154;
razn_w_mem[11311] = 154;
razn_w_mem[11312] = 154;
razn_w_mem[11313] = 154;
razn_w_mem[11314] = 154;
razn_w_mem[11315] = 154;
razn_w_mem[11316] = 154;
razn_w_mem[11317] = 154;
razn_w_mem[11318] = 154;
razn_w_mem[11319] = 154;
razn_w_mem[11320] = 154;
razn_w_mem[11321] = 154;
razn_w_mem[11322] = 154;
razn_w_mem[11323] = 154;
razn_w_mem[11324] = 154;
razn_w_mem[11325] = 154;
razn_w_mem[11326] = 154;
razn_w_mem[11327] = 154;
razn_w_mem[11328] = 154;
razn_w_mem[11329] = 154;
razn_w_mem[11330] = 154;
razn_w_mem[11331] = 154;
razn_w_mem[11332] = 154;
razn_w_mem[11333] = 154;
razn_w_mem[11334] = 154;
razn_w_mem[11335] = 154;
razn_w_mem[11336] = 154;
razn_w_mem[11337] = 154;
razn_w_mem[11338] = 154;
razn_w_mem[11339] = 154;
razn_w_mem[11340] = 154;
razn_w_mem[11341] = 154;
razn_w_mem[11342] = 154;
razn_w_mem[11343] = 154;
razn_w_mem[11344] = 154;
razn_w_mem[11345] = 154;
razn_w_mem[11346] = 154;
razn_w_mem[11347] = 154;
razn_w_mem[11348] = 154;
razn_w_mem[11349] = 154;
razn_w_mem[11350] = 154;
razn_w_mem[11351] = 154;
razn_w_mem[11352] = 154;
razn_w_mem[11353] = 154;
razn_w_mem[11354] = 154;
razn_w_mem[11355] = 154;
razn_w_mem[11356] = 154;
razn_w_mem[11357] = 154;
razn_w_mem[11358] = 154;
razn_w_mem[11359] = 154;
razn_w_mem[11360] = 154;
razn_w_mem[11361] = 154;
razn_w_mem[11362] = 154;
razn_w_mem[11363] = 154;
razn_w_mem[11364] = 154;
razn_w_mem[11365] = 154;
razn_w_mem[11366] = 154;
razn_w_mem[11367] = 154;
razn_w_mem[11368] = 154;
razn_w_mem[11369] = 154;
razn_w_mem[11370] = 154;
razn_w_mem[11371] = 154;
razn_w_mem[11372] = 154;
razn_w_mem[11373] = 154;
razn_w_mem[11374] = 154;
razn_w_mem[11375] = 154;
razn_w_mem[11376] = 154;
razn_w_mem[11377] = 154;
razn_w_mem[11378] = 154;
razn_w_mem[11379] = 154;
razn_w_mem[11380] = 154;
razn_w_mem[11381] = 154;
razn_w_mem[11382] = 154;
razn_w_mem[11383] = 154;
razn_w_mem[11384] = 154;
razn_w_mem[11385] = 154;
razn_w_mem[11386] = 154;
razn_w_mem[11387] = 154;
razn_w_mem[11388] = 154;
razn_w_mem[11389] = 154;
razn_w_mem[11390] = 154;
razn_w_mem[11391] = 154;
razn_w_mem[11392] = 124;
razn_w_mem[11393] = 124;
razn_w_mem[11394] = 124;
razn_w_mem[11395] = 124;
razn_w_mem[11396] = 124;
razn_w_mem[11397] = 124;
razn_w_mem[11398] = 124;
razn_w_mem[11399] = 124;
razn_w_mem[11400] = 124;
razn_w_mem[11401] = 124;
razn_w_mem[11402] = 124;
razn_w_mem[11403] = 124;
razn_w_mem[11404] = 124;
razn_w_mem[11405] = 124;
razn_w_mem[11406] = 124;
razn_w_mem[11407] = 124;
razn_w_mem[11408] = 124;
razn_w_mem[11409] = 124;
razn_w_mem[11410] = 124;
razn_w_mem[11411] = 124;
razn_w_mem[11412] = 124;
razn_w_mem[11413] = 124;
razn_w_mem[11414] = 124;
razn_w_mem[11415] = 124;
razn_w_mem[11416] = 124;
razn_w_mem[11417] = 124;
razn_w_mem[11418] = 124;
razn_w_mem[11419] = 124;
razn_w_mem[11420] = 124;
razn_w_mem[11421] = 124;
razn_w_mem[11422] = 124;
razn_w_mem[11423] = 124;
razn_w_mem[11424] = 124;
razn_w_mem[11425] = 124;
razn_w_mem[11426] = 124;
razn_w_mem[11427] = 124;
razn_w_mem[11428] = 124;
razn_w_mem[11429] = 124;
razn_w_mem[11430] = 124;
razn_w_mem[11431] = 124;
razn_w_mem[11432] = 124;
razn_w_mem[11433] = 124;
razn_w_mem[11434] = 124;
razn_w_mem[11435] = 124;
razn_w_mem[11436] = 124;
razn_w_mem[11437] = 124;
razn_w_mem[11438] = 124;
razn_w_mem[11439] = 124;
razn_w_mem[11440] = 124;
razn_w_mem[11441] = 124;
razn_w_mem[11442] = 124;
razn_w_mem[11443] = 124;
razn_w_mem[11444] = 124;
razn_w_mem[11445] = 124;
razn_w_mem[11446] = 124;
razn_w_mem[11447] = 124;
razn_w_mem[11448] = 124;
razn_w_mem[11449] = 124;
razn_w_mem[11450] = 124;
razn_w_mem[11451] = 124;
razn_w_mem[11452] = 124;
razn_w_mem[11453] = 124;
razn_w_mem[11454] = 124;
razn_w_mem[11455] = 124;
razn_w_mem[11456] = 124;
razn_w_mem[11457] = 124;
razn_w_mem[11458] = 124;
razn_w_mem[11459] = 124;
razn_w_mem[11460] = 124;
razn_w_mem[11461] = 124;
razn_w_mem[11462] = 124;
razn_w_mem[11463] = 124;
razn_w_mem[11464] = 124;
razn_w_mem[11465] = 124;
razn_w_mem[11466] = 124;
razn_w_mem[11467] = 124;
razn_w_mem[11468] = 124;
razn_w_mem[11469] = 124;
razn_w_mem[11470] = 124;
razn_w_mem[11471] = 124;
razn_w_mem[11472] = 124;
razn_w_mem[11473] = 124;
razn_w_mem[11474] = 124;
razn_w_mem[11475] = 124;
razn_w_mem[11476] = 124;
razn_w_mem[11477] = 124;
razn_w_mem[11478] = 124;
razn_w_mem[11479] = 124;
razn_w_mem[11480] = 124;
razn_w_mem[11481] = 124;
razn_w_mem[11482] = 124;
razn_w_mem[11483] = 124;
razn_w_mem[11484] = 124;
razn_w_mem[11485] = 124;
razn_w_mem[11486] = 124;
razn_w_mem[11487] = 124;
razn_w_mem[11488] = 124;
razn_w_mem[11489] = 124;
razn_w_mem[11490] = 124;
razn_w_mem[11491] = 124;
razn_w_mem[11492] = 124;
razn_w_mem[11493] = 124;
razn_w_mem[11494] = 124;
razn_w_mem[11495] = 124;
razn_w_mem[11496] = 124;
razn_w_mem[11497] = 124;
razn_w_mem[11498] = 124;
razn_w_mem[11499] = 124;
razn_w_mem[11500] = 124;
razn_w_mem[11501] = 124;
razn_w_mem[11502] = 124;
razn_w_mem[11503] = 124;
razn_w_mem[11504] = 124;
razn_w_mem[11505] = 124;
razn_w_mem[11506] = 124;
razn_w_mem[11507] = 124;
razn_w_mem[11508] = 124;
razn_w_mem[11509] = 124;
razn_w_mem[11510] = 124;
razn_w_mem[11511] = 124;
razn_w_mem[11512] = 124;
razn_w_mem[11513] = 124;
razn_w_mem[11514] = 124;
razn_w_mem[11515] = 124;
razn_w_mem[11516] = 124;
razn_w_mem[11517] = 124;
razn_w_mem[11518] = 124;
razn_w_mem[11519] = 124;
razn_w_mem[11520] = 94;
razn_w_mem[11521] = 94;
razn_w_mem[11522] = 94;
razn_w_mem[11523] = 94;
razn_w_mem[11524] = 94;
razn_w_mem[11525] = 94;
razn_w_mem[11526] = 94;
razn_w_mem[11527] = 94;
razn_w_mem[11528] = 94;
razn_w_mem[11529] = 94;
razn_w_mem[11530] = 94;
razn_w_mem[11531] = 94;
razn_w_mem[11532] = 94;
razn_w_mem[11533] = 94;
razn_w_mem[11534] = 94;
razn_w_mem[11535] = 94;
razn_w_mem[11536] = 94;
razn_w_mem[11537] = 94;
razn_w_mem[11538] = 94;
razn_w_mem[11539] = 94;
razn_w_mem[11540] = 94;
razn_w_mem[11541] = 94;
razn_w_mem[11542] = 94;
razn_w_mem[11543] = 94;
razn_w_mem[11544] = 94;
razn_w_mem[11545] = 94;
razn_w_mem[11546] = 94;
razn_w_mem[11547] = 94;
razn_w_mem[11548] = 94;
razn_w_mem[11549] = 94;
razn_w_mem[11550] = 94;
razn_w_mem[11551] = 94;
razn_w_mem[11552] = 94;
razn_w_mem[11553] = 94;
razn_w_mem[11554] = 94;
razn_w_mem[11555] = 94;
razn_w_mem[11556] = 94;
razn_w_mem[11557] = 94;
razn_w_mem[11558] = 94;
razn_w_mem[11559] = 94;
razn_w_mem[11560] = 94;
razn_w_mem[11561] = 94;
razn_w_mem[11562] = 94;
razn_w_mem[11563] = 94;
razn_w_mem[11564] = 94;
razn_w_mem[11565] = 94;
razn_w_mem[11566] = 94;
razn_w_mem[11567] = 94;
razn_w_mem[11568] = 94;
razn_w_mem[11569] = 94;
razn_w_mem[11570] = 94;
razn_w_mem[11571] = 94;
razn_w_mem[11572] = 94;
razn_w_mem[11573] = 94;
razn_w_mem[11574] = 94;
razn_w_mem[11575] = 94;
razn_w_mem[11576] = 94;
razn_w_mem[11577] = 94;
razn_w_mem[11578] = 94;
razn_w_mem[11579] = 94;
razn_w_mem[11580] = 94;
razn_w_mem[11581] = 94;
razn_w_mem[11582] = 94;
razn_w_mem[11583] = 94;
razn_w_mem[11584] = 94;
razn_w_mem[11585] = 94;
razn_w_mem[11586] = 94;
razn_w_mem[11587] = 94;
razn_w_mem[11588] = 94;
razn_w_mem[11589] = 94;
razn_w_mem[11590] = 94;
razn_w_mem[11591] = 94;
razn_w_mem[11592] = 94;
razn_w_mem[11593] = 94;
razn_w_mem[11594] = 94;
razn_w_mem[11595] = 94;
razn_w_mem[11596] = 94;
razn_w_mem[11597] = 94;
razn_w_mem[11598] = 94;
razn_w_mem[11599] = 94;
razn_w_mem[11600] = 94;
razn_w_mem[11601] = 94;
razn_w_mem[11602] = 94;
razn_w_mem[11603] = 94;
razn_w_mem[11604] = 94;
razn_w_mem[11605] = 94;
razn_w_mem[11606] = 94;
razn_w_mem[11607] = 94;
razn_w_mem[11608] = 94;
razn_w_mem[11609] = 94;
razn_w_mem[11610] = 94;
razn_w_mem[11611] = 94;
razn_w_mem[11612] = 94;
razn_w_mem[11613] = 94;
razn_w_mem[11614] = 94;
razn_w_mem[11615] = 94;
razn_w_mem[11616] = 94;
razn_w_mem[11617] = 94;
razn_w_mem[11618] = 94;
razn_w_mem[11619] = 94;
razn_w_mem[11620] = 94;
razn_w_mem[11621] = 94;
razn_w_mem[11622] = 94;
razn_w_mem[11623] = 94;
razn_w_mem[11624] = 94;
razn_w_mem[11625] = 94;
razn_w_mem[11626] = 94;
razn_w_mem[11627] = 94;
razn_w_mem[11628] = 94;
razn_w_mem[11629] = 94;
razn_w_mem[11630] = 94;
razn_w_mem[11631] = 94;
razn_w_mem[11632] = 94;
razn_w_mem[11633] = 94;
razn_w_mem[11634] = 94;
razn_w_mem[11635] = 94;
razn_w_mem[11636] = 94;
razn_w_mem[11637] = 94;
razn_w_mem[11638] = 94;
razn_w_mem[11639] = 94;
razn_w_mem[11640] = 94;
razn_w_mem[11641] = 94;
razn_w_mem[11642] = 94;
razn_w_mem[11643] = 94;
razn_w_mem[11644] = 94;
razn_w_mem[11645] = 94;
razn_w_mem[11646] = 94;
razn_w_mem[11647] = 94;
razn_w_mem[11648] = 64;
razn_w_mem[11649] = 64;
razn_w_mem[11650] = 64;
razn_w_mem[11651] = 64;
razn_w_mem[11652] = 64;
razn_w_mem[11653] = 64;
razn_w_mem[11654] = 64;
razn_w_mem[11655] = 64;
razn_w_mem[11656] = 64;
razn_w_mem[11657] = 64;
razn_w_mem[11658] = 64;
razn_w_mem[11659] = 64;
razn_w_mem[11660] = 64;
razn_w_mem[11661] = 64;
razn_w_mem[11662] = 64;
razn_w_mem[11663] = 64;
razn_w_mem[11664] = 64;
razn_w_mem[11665] = 64;
razn_w_mem[11666] = 64;
razn_w_mem[11667] = 64;
razn_w_mem[11668] = 64;
razn_w_mem[11669] = 64;
razn_w_mem[11670] = 64;
razn_w_mem[11671] = 64;
razn_w_mem[11672] = 64;
razn_w_mem[11673] = 64;
razn_w_mem[11674] = 64;
razn_w_mem[11675] = 64;
razn_w_mem[11676] = 64;
razn_w_mem[11677] = 64;
razn_w_mem[11678] = 64;
razn_w_mem[11679] = 64;
razn_w_mem[11680] = 64;
razn_w_mem[11681] = 64;
razn_w_mem[11682] = 64;
razn_w_mem[11683] = 64;
razn_w_mem[11684] = 64;
razn_w_mem[11685] = 64;
razn_w_mem[11686] = 64;
razn_w_mem[11687] = 64;
razn_w_mem[11688] = 64;
razn_w_mem[11689] = 64;
razn_w_mem[11690] = 64;
razn_w_mem[11691] = 64;
razn_w_mem[11692] = 64;
razn_w_mem[11693] = 64;
razn_w_mem[11694] = 64;
razn_w_mem[11695] = 64;
razn_w_mem[11696] = 64;
razn_w_mem[11697] = 64;
razn_w_mem[11698] = 64;
razn_w_mem[11699] = 64;
razn_w_mem[11700] = 64;
razn_w_mem[11701] = 64;
razn_w_mem[11702] = 64;
razn_w_mem[11703] = 64;
razn_w_mem[11704] = 64;
razn_w_mem[11705] = 64;
razn_w_mem[11706] = 64;
razn_w_mem[11707] = 64;
razn_w_mem[11708] = 64;
razn_w_mem[11709] = 64;
razn_w_mem[11710] = 64;
razn_w_mem[11711] = 64;
razn_w_mem[11712] = 64;
razn_w_mem[11713] = 64;
razn_w_mem[11714] = 64;
razn_w_mem[11715] = 64;
razn_w_mem[11716] = 64;
razn_w_mem[11717] = 64;
razn_w_mem[11718] = 64;
razn_w_mem[11719] = 64;
razn_w_mem[11720] = 64;
razn_w_mem[11721] = 64;
razn_w_mem[11722] = 64;
razn_w_mem[11723] = 64;
razn_w_mem[11724] = 64;
razn_w_mem[11725] = 64;
razn_w_mem[11726] = 64;
razn_w_mem[11727] = 64;
razn_w_mem[11728] = 64;
razn_w_mem[11729] = 64;
razn_w_mem[11730] = 64;
razn_w_mem[11731] = 64;
razn_w_mem[11732] = 64;
razn_w_mem[11733] = 64;
razn_w_mem[11734] = 64;
razn_w_mem[11735] = 64;
razn_w_mem[11736] = 64;
razn_w_mem[11737] = 64;
razn_w_mem[11738] = 64;
razn_w_mem[11739] = 64;
razn_w_mem[11740] = 64;
razn_w_mem[11741] = 64;
razn_w_mem[11742] = 64;
razn_w_mem[11743] = 64;
razn_w_mem[11744] = 64;
razn_w_mem[11745] = 64;
razn_w_mem[11746] = 64;
razn_w_mem[11747] = 64;
razn_w_mem[11748] = 64;
razn_w_mem[11749] = 64;
razn_w_mem[11750] = 64;
razn_w_mem[11751] = 64;
razn_w_mem[11752] = 64;
razn_w_mem[11753] = 64;
razn_w_mem[11754] = 64;
razn_w_mem[11755] = 64;
razn_w_mem[11756] = 64;
razn_w_mem[11757] = 64;
razn_w_mem[11758] = 64;
razn_w_mem[11759] = 64;
razn_w_mem[11760] = 64;
razn_w_mem[11761] = 64;
razn_w_mem[11762] = 64;
razn_w_mem[11763] = 64;
razn_w_mem[11764] = 64;
razn_w_mem[11765] = 64;
razn_w_mem[11766] = 64;
razn_w_mem[11767] = 64;
razn_w_mem[11768] = 64;
razn_w_mem[11769] = 64;
razn_w_mem[11770] = 64;
razn_w_mem[11771] = 64;
razn_w_mem[11772] = 64;
razn_w_mem[11773] = 64;
razn_w_mem[11774] = 64;
razn_w_mem[11775] = 64;
razn_w_mem[11776] = 34;
razn_w_mem[11777] = 34;
razn_w_mem[11778] = 34;
razn_w_mem[11779] = 34;
razn_w_mem[11780] = 34;
razn_w_mem[11781] = 34;
razn_w_mem[11782] = 34;
razn_w_mem[11783] = 34;
razn_w_mem[11784] = 34;
razn_w_mem[11785] = 34;
razn_w_mem[11786] = 34;
razn_w_mem[11787] = 34;
razn_w_mem[11788] = 34;
razn_w_mem[11789] = 34;
razn_w_mem[11790] = 34;
razn_w_mem[11791] = 34;
razn_w_mem[11792] = 34;
razn_w_mem[11793] = 34;
razn_w_mem[11794] = 34;
razn_w_mem[11795] = 34;
razn_w_mem[11796] = 34;
razn_w_mem[11797] = 34;
razn_w_mem[11798] = 34;
razn_w_mem[11799] = 34;
razn_w_mem[11800] = 34;
razn_w_mem[11801] = 34;
razn_w_mem[11802] = 34;
razn_w_mem[11803] = 34;
razn_w_mem[11804] = 34;
razn_w_mem[11805] = 34;
razn_w_mem[11806] = 34;
razn_w_mem[11807] = 34;
razn_w_mem[11808] = 34;
razn_w_mem[11809] = 34;
razn_w_mem[11810] = 34;
razn_w_mem[11811] = 34;
razn_w_mem[11812] = 34;
razn_w_mem[11813] = 34;
razn_w_mem[11814] = 34;
razn_w_mem[11815] = 34;
razn_w_mem[11816] = 34;
razn_w_mem[11817] = 34;
razn_w_mem[11818] = 34;
razn_w_mem[11819] = 34;
razn_w_mem[11820] = 34;
razn_w_mem[11821] = 34;
razn_w_mem[11822] = 34;
razn_w_mem[11823] = 34;
razn_w_mem[11824] = 34;
razn_w_mem[11825] = 34;
razn_w_mem[11826] = 34;
razn_w_mem[11827] = 34;
razn_w_mem[11828] = 34;
razn_w_mem[11829] = 34;
razn_w_mem[11830] = 34;
razn_w_mem[11831] = 34;
razn_w_mem[11832] = 34;
razn_w_mem[11833] = 34;
razn_w_mem[11834] = 34;
razn_w_mem[11835] = 34;
razn_w_mem[11836] = 34;
razn_w_mem[11837] = 34;
razn_w_mem[11838] = 34;
razn_w_mem[11839] = 34;
razn_w_mem[11840] = 34;
razn_w_mem[11841] = 34;
razn_w_mem[11842] = 34;
razn_w_mem[11843] = 34;
razn_w_mem[11844] = 34;
razn_w_mem[11845] = 34;
razn_w_mem[11846] = 34;
razn_w_mem[11847] = 34;
razn_w_mem[11848] = 34;
razn_w_mem[11849] = 34;
razn_w_mem[11850] = 34;
razn_w_mem[11851] = 34;
razn_w_mem[11852] = 34;
razn_w_mem[11853] = 34;
razn_w_mem[11854] = 34;
razn_w_mem[11855] = 34;
razn_w_mem[11856] = 34;
razn_w_mem[11857] = 34;
razn_w_mem[11858] = 34;
razn_w_mem[11859] = 34;
razn_w_mem[11860] = 34;
razn_w_mem[11861] = 34;
razn_w_mem[11862] = 34;
razn_w_mem[11863] = 34;
razn_w_mem[11864] = 34;
razn_w_mem[11865] = 34;
razn_w_mem[11866] = 34;
razn_w_mem[11867] = 34;
razn_w_mem[11868] = 34;
razn_w_mem[11869] = 34;
razn_w_mem[11870] = 34;
razn_w_mem[11871] = 34;
razn_w_mem[11872] = 34;
razn_w_mem[11873] = 34;
razn_w_mem[11874] = 34;
razn_w_mem[11875] = 34;
razn_w_mem[11876] = 34;
razn_w_mem[11877] = 34;
razn_w_mem[11878] = 34;
razn_w_mem[11879] = 34;
razn_w_mem[11880] = 34;
razn_w_mem[11881] = 34;
razn_w_mem[11882] = 34;
razn_w_mem[11883] = 34;
razn_w_mem[11884] = 34;
razn_w_mem[11885] = 34;
razn_w_mem[11886] = 34;
razn_w_mem[11887] = 34;
razn_w_mem[11888] = 34;
razn_w_mem[11889] = 34;
razn_w_mem[11890] = 34;
razn_w_mem[11891] = 34;
razn_w_mem[11892] = 34;
razn_w_mem[11893] = 34;
razn_w_mem[11894] = 34;
razn_w_mem[11895] = 34;
razn_w_mem[11896] = 34;
razn_w_mem[11897] = 34;
razn_w_mem[11898] = 34;
razn_w_mem[11899] = 34;
razn_w_mem[11900] = 34;
razn_w_mem[11901] = 34;
razn_w_mem[11902] = 34;
razn_w_mem[11903] = 34;
razn_w_mem[11904] = 4;
razn_w_mem[11905] = 4;
razn_w_mem[11906] = 4;
razn_w_mem[11907] = 4;
razn_w_mem[11908] = 4;
razn_w_mem[11909] = 4;
razn_w_mem[11910] = 4;
razn_w_mem[11911] = 4;
razn_w_mem[11912] = 4;
razn_w_mem[11913] = 4;
razn_w_mem[11914] = 4;
razn_w_mem[11915] = 4;
razn_w_mem[11916] = 4;
razn_w_mem[11917] = 4;
razn_w_mem[11918] = 4;
razn_w_mem[11919] = 4;
razn_w_mem[11920] = 4;
razn_w_mem[11921] = 4;
razn_w_mem[11922] = 4;
razn_w_mem[11923] = 4;
razn_w_mem[11924] = 4;
razn_w_mem[11925] = 4;
razn_w_mem[11926] = 4;
razn_w_mem[11927] = 4;
razn_w_mem[11928] = 4;
razn_w_mem[11929] = 4;
razn_w_mem[11930] = 4;
razn_w_mem[11931] = 4;
razn_w_mem[11932] = 4;
razn_w_mem[11933] = 4;
razn_w_mem[11934] = 4;
razn_w_mem[11935] = 4;
razn_w_mem[11936] = 4;
razn_w_mem[11937] = 4;
razn_w_mem[11938] = 4;
razn_w_mem[11939] = 4;
razn_w_mem[11940] = 4;
razn_w_mem[11941] = 4;
razn_w_mem[11942] = 4;
razn_w_mem[11943] = 4;
razn_w_mem[11944] = 4;
razn_w_mem[11945] = 4;
razn_w_mem[11946] = 4;
razn_w_mem[11947] = 4;
razn_w_mem[11948] = 4;
razn_w_mem[11949] = 4;
razn_w_mem[11950] = 4;
razn_w_mem[11951] = 4;
razn_w_mem[11952] = 4;
razn_w_mem[11953] = 4;
razn_w_mem[11954] = 4;
razn_w_mem[11955] = 4;
razn_w_mem[11956] = 4;
razn_w_mem[11957] = 4;
razn_w_mem[11958] = 4;
razn_w_mem[11959] = 4;
razn_w_mem[11960] = 4;
razn_w_mem[11961] = 4;
razn_w_mem[11962] = 4;
razn_w_mem[11963] = 4;
razn_w_mem[11964] = 4;
razn_w_mem[11965] = 4;
razn_w_mem[11966] = 4;
razn_w_mem[11967] = 4;
razn_w_mem[11968] = 4;
razn_w_mem[11969] = 4;
razn_w_mem[11970] = 4;
razn_w_mem[11971] = 4;
razn_w_mem[11972] = 4;
razn_w_mem[11973] = 4;
razn_w_mem[11974] = 4;
razn_w_mem[11975] = 4;
razn_w_mem[11976] = 4;
razn_w_mem[11977] = 4;
razn_w_mem[11978] = 4;
razn_w_mem[11979] = 4;
razn_w_mem[11980] = 4;
razn_w_mem[11981] = 4;
razn_w_mem[11982] = 4;
razn_w_mem[11983] = 4;
razn_w_mem[11984] = 4;
razn_w_mem[11985] = 4;
razn_w_mem[11986] = 4;
razn_w_mem[11987] = 4;
razn_w_mem[11988] = 4;
razn_w_mem[11989] = 4;
razn_w_mem[11990] = 4;
razn_w_mem[11991] = 4;
razn_w_mem[11992] = 4;
razn_w_mem[11993] = 4;
razn_w_mem[11994] = 4;
razn_w_mem[11995] = 4;
razn_w_mem[11996] = 4;
razn_w_mem[11997] = 4;
razn_w_mem[11998] = 4;
razn_w_mem[11999] = 4;
razn_w_mem[12000] = 4;
razn_w_mem[12001] = 4;
razn_w_mem[12002] = 4;
razn_w_mem[12003] = 4;
razn_w_mem[12004] = 4;
razn_w_mem[12005] = 4;
razn_w_mem[12006] = 4;
razn_w_mem[12007] = 4;
razn_w_mem[12008] = 4;
razn_w_mem[12009] = 4;
razn_w_mem[12010] = 4;
razn_w_mem[12011] = 4;
razn_w_mem[12012] = 4;
razn_w_mem[12013] = 4;
razn_w_mem[12014] = 4;
razn_w_mem[12015] = 4;
razn_w_mem[12016] = 4;
razn_w_mem[12017] = 4;
razn_w_mem[12018] = 4;
razn_w_mem[12019] = 4;
razn_w_mem[12020] = 4;
razn_w_mem[12021] = 4;
razn_w_mem[12022] = 4;
razn_w_mem[12023] = 4;
razn_w_mem[12024] = 4;
razn_w_mem[12025] = 4;
razn_w_mem[12026] = 4;
razn_w_mem[12027] = 4;
razn_w_mem[12028] = 4;
razn_w_mem[12029] = 4;
razn_w_mem[12030] = 4;
razn_w_mem[12031] = 4;
razn_w_mem[12032] = 228;
razn_w_mem[12033] = 228;
razn_w_mem[12034] = 228;
razn_w_mem[12035] = 228;
razn_w_mem[12036] = 228;
razn_w_mem[12037] = 228;
razn_w_mem[12038] = 228;
razn_w_mem[12039] = 228;
razn_w_mem[12040] = 228;
razn_w_mem[12041] = 228;
razn_w_mem[12042] = 228;
razn_w_mem[12043] = 228;
razn_w_mem[12044] = 228;
razn_w_mem[12045] = 228;
razn_w_mem[12046] = 228;
razn_w_mem[12047] = 228;
razn_w_mem[12048] = 228;
razn_w_mem[12049] = 228;
razn_w_mem[12050] = 228;
razn_w_mem[12051] = 228;
razn_w_mem[12052] = 228;
razn_w_mem[12053] = 228;
razn_w_mem[12054] = 228;
razn_w_mem[12055] = 228;
razn_w_mem[12056] = 228;
razn_w_mem[12057] = 228;
razn_w_mem[12058] = 228;
razn_w_mem[12059] = 228;
razn_w_mem[12060] = 228;
razn_w_mem[12061] = 228;
razn_w_mem[12062] = 228;
razn_w_mem[12063] = 228;
razn_w_mem[12064] = 228;
razn_w_mem[12065] = 228;
razn_w_mem[12066] = 228;
razn_w_mem[12067] = 228;
razn_w_mem[12068] = 228;
razn_w_mem[12069] = 228;
razn_w_mem[12070] = 228;
razn_w_mem[12071] = 228;
razn_w_mem[12072] = 228;
razn_w_mem[12073] = 228;
razn_w_mem[12074] = 228;
razn_w_mem[12075] = 228;
razn_w_mem[12076] = 228;
razn_w_mem[12077] = 228;
razn_w_mem[12078] = 228;
razn_w_mem[12079] = 228;
razn_w_mem[12080] = 228;
razn_w_mem[12081] = 228;
razn_w_mem[12082] = 228;
razn_w_mem[12083] = 228;
razn_w_mem[12084] = 228;
razn_w_mem[12085] = 228;
razn_w_mem[12086] = 228;
razn_w_mem[12087] = 228;
razn_w_mem[12088] = 228;
razn_w_mem[12089] = 228;
razn_w_mem[12090] = 228;
razn_w_mem[12091] = 228;
razn_w_mem[12092] = 228;
razn_w_mem[12093] = 228;
razn_w_mem[12094] = 228;
razn_w_mem[12095] = 228;
razn_w_mem[12096] = 228;
razn_w_mem[12097] = 228;
razn_w_mem[12098] = 228;
razn_w_mem[12099] = 228;
razn_w_mem[12100] = 228;
razn_w_mem[12101] = 228;
razn_w_mem[12102] = 228;
razn_w_mem[12103] = 228;
razn_w_mem[12104] = 228;
razn_w_mem[12105] = 228;
razn_w_mem[12106] = 228;
razn_w_mem[12107] = 228;
razn_w_mem[12108] = 228;
razn_w_mem[12109] = 228;
razn_w_mem[12110] = 228;
razn_w_mem[12111] = 228;
razn_w_mem[12112] = 228;
razn_w_mem[12113] = 228;
razn_w_mem[12114] = 228;
razn_w_mem[12115] = 228;
razn_w_mem[12116] = 228;
razn_w_mem[12117] = 228;
razn_w_mem[12118] = 228;
razn_w_mem[12119] = 228;
razn_w_mem[12120] = 228;
razn_w_mem[12121] = 228;
razn_w_mem[12122] = 228;
razn_w_mem[12123] = 228;
razn_w_mem[12124] = 228;
razn_w_mem[12125] = 228;
razn_w_mem[12126] = 228;
razn_w_mem[12127] = 228;
razn_w_mem[12128] = 228;
razn_w_mem[12129] = 228;
razn_w_mem[12130] = 228;
razn_w_mem[12131] = 228;
razn_w_mem[12132] = 228;
razn_w_mem[12133] = 228;
razn_w_mem[12134] = 228;
razn_w_mem[12135] = 228;
razn_w_mem[12136] = 228;
razn_w_mem[12137] = 228;
razn_w_mem[12138] = 228;
razn_w_mem[12139] = 228;
razn_w_mem[12140] = 228;
razn_w_mem[12141] = 228;
razn_w_mem[12142] = 228;
razn_w_mem[12143] = 228;
razn_w_mem[12144] = 228;
razn_w_mem[12145] = 228;
razn_w_mem[12146] = 228;
razn_w_mem[12147] = 228;
razn_w_mem[12148] = 228;
razn_w_mem[12149] = 228;
razn_w_mem[12150] = 228;
razn_w_mem[12151] = 228;
razn_w_mem[12152] = 228;
razn_w_mem[12153] = 228;
razn_w_mem[12154] = 228;
razn_w_mem[12155] = 228;
razn_w_mem[12156] = 228;
razn_w_mem[12157] = 228;
razn_w_mem[12158] = 228;
razn_w_mem[12159] = 228;
razn_w_mem[12160] = 198;
razn_w_mem[12161] = 198;
razn_w_mem[12162] = 198;
razn_w_mem[12163] = 198;
razn_w_mem[12164] = 198;
razn_w_mem[12165] = 198;
razn_w_mem[12166] = 198;
razn_w_mem[12167] = 198;
razn_w_mem[12168] = 198;
razn_w_mem[12169] = 198;
razn_w_mem[12170] = 198;
razn_w_mem[12171] = 198;
razn_w_mem[12172] = 198;
razn_w_mem[12173] = 198;
razn_w_mem[12174] = 198;
razn_w_mem[12175] = 198;
razn_w_mem[12176] = 198;
razn_w_mem[12177] = 198;
razn_w_mem[12178] = 198;
razn_w_mem[12179] = 198;
razn_w_mem[12180] = 198;
razn_w_mem[12181] = 198;
razn_w_mem[12182] = 198;
razn_w_mem[12183] = 198;
razn_w_mem[12184] = 198;
razn_w_mem[12185] = 198;
razn_w_mem[12186] = 198;
razn_w_mem[12187] = 198;
razn_w_mem[12188] = 198;
razn_w_mem[12189] = 198;
razn_w_mem[12190] = 198;
razn_w_mem[12191] = 198;
razn_w_mem[12192] = 198;
razn_w_mem[12193] = 198;
razn_w_mem[12194] = 198;
razn_w_mem[12195] = 198;
razn_w_mem[12196] = 198;
razn_w_mem[12197] = 198;
razn_w_mem[12198] = 198;
razn_w_mem[12199] = 198;
razn_w_mem[12200] = 198;
razn_w_mem[12201] = 198;
razn_w_mem[12202] = 198;
razn_w_mem[12203] = 198;
razn_w_mem[12204] = 198;
razn_w_mem[12205] = 198;
razn_w_mem[12206] = 198;
razn_w_mem[12207] = 198;
razn_w_mem[12208] = 198;
razn_w_mem[12209] = 198;
razn_w_mem[12210] = 198;
razn_w_mem[12211] = 198;
razn_w_mem[12212] = 198;
razn_w_mem[12213] = 198;
razn_w_mem[12214] = 198;
razn_w_mem[12215] = 198;
razn_w_mem[12216] = 198;
razn_w_mem[12217] = 198;
razn_w_mem[12218] = 198;
razn_w_mem[12219] = 198;
razn_w_mem[12220] = 198;
razn_w_mem[12221] = 198;
razn_w_mem[12222] = 198;
razn_w_mem[12223] = 198;
razn_w_mem[12224] = 198;
razn_w_mem[12225] = 198;
razn_w_mem[12226] = 198;
razn_w_mem[12227] = 198;
razn_w_mem[12228] = 198;
razn_w_mem[12229] = 198;
razn_w_mem[12230] = 198;
razn_w_mem[12231] = 198;
razn_w_mem[12232] = 198;
razn_w_mem[12233] = 198;
razn_w_mem[12234] = 198;
razn_w_mem[12235] = 198;
razn_w_mem[12236] = 198;
razn_w_mem[12237] = 198;
razn_w_mem[12238] = 198;
razn_w_mem[12239] = 198;
razn_w_mem[12240] = 198;
razn_w_mem[12241] = 198;
razn_w_mem[12242] = 198;
razn_w_mem[12243] = 198;
razn_w_mem[12244] = 198;
razn_w_mem[12245] = 198;
razn_w_mem[12246] = 198;
razn_w_mem[12247] = 198;
razn_w_mem[12248] = 198;
razn_w_mem[12249] = 198;
razn_w_mem[12250] = 198;
razn_w_mem[12251] = 198;
razn_w_mem[12252] = 198;
razn_w_mem[12253] = 198;
razn_w_mem[12254] = 198;
razn_w_mem[12255] = 198;
razn_w_mem[12256] = 198;
razn_w_mem[12257] = 198;
razn_w_mem[12258] = 198;
razn_w_mem[12259] = 198;
razn_w_mem[12260] = 198;
razn_w_mem[12261] = 198;
razn_w_mem[12262] = 198;
razn_w_mem[12263] = 198;
razn_w_mem[12264] = 198;
razn_w_mem[12265] = 198;
razn_w_mem[12266] = 198;
razn_w_mem[12267] = 198;
razn_w_mem[12268] = 198;
razn_w_mem[12269] = 198;
razn_w_mem[12270] = 198;
razn_w_mem[12271] = 198;
razn_w_mem[12272] = 198;
razn_w_mem[12273] = 198;
razn_w_mem[12274] = 198;
razn_w_mem[12275] = 198;
razn_w_mem[12276] = 198;
razn_w_mem[12277] = 198;
razn_w_mem[12278] = 198;
razn_w_mem[12279] = 198;
razn_w_mem[12280] = 198;
razn_w_mem[12281] = 198;
razn_w_mem[12282] = 198;
razn_w_mem[12283] = 198;
razn_w_mem[12284] = 198;
razn_w_mem[12285] = 198;
razn_w_mem[12286] = 198;
razn_w_mem[12287] = 198;
razn_w_mem[12288] = 168;
razn_w_mem[12289] = 168;
razn_w_mem[12290] = 168;
razn_w_mem[12291] = 168;
razn_w_mem[12292] = 168;
razn_w_mem[12293] = 168;
razn_w_mem[12294] = 168;
razn_w_mem[12295] = 168;
razn_w_mem[12296] = 168;
razn_w_mem[12297] = 168;
razn_w_mem[12298] = 168;
razn_w_mem[12299] = 168;
razn_w_mem[12300] = 168;
razn_w_mem[12301] = 168;
razn_w_mem[12302] = 168;
razn_w_mem[12303] = 168;
razn_w_mem[12304] = 168;
razn_w_mem[12305] = 168;
razn_w_mem[12306] = 168;
razn_w_mem[12307] = 168;
razn_w_mem[12308] = 168;
razn_w_mem[12309] = 168;
razn_w_mem[12310] = 168;
razn_w_mem[12311] = 168;
razn_w_mem[12312] = 168;
razn_w_mem[12313] = 168;
razn_w_mem[12314] = 168;
razn_w_mem[12315] = 168;
razn_w_mem[12316] = 168;
razn_w_mem[12317] = 168;
razn_w_mem[12318] = 168;
razn_w_mem[12319] = 168;
razn_w_mem[12320] = 168;
razn_w_mem[12321] = 168;
razn_w_mem[12322] = 168;
razn_w_mem[12323] = 168;
razn_w_mem[12324] = 168;
razn_w_mem[12325] = 168;
razn_w_mem[12326] = 168;
razn_w_mem[12327] = 168;
razn_w_mem[12328] = 168;
razn_w_mem[12329] = 168;
razn_w_mem[12330] = 168;
razn_w_mem[12331] = 168;
razn_w_mem[12332] = 168;
razn_w_mem[12333] = 168;
razn_w_mem[12334] = 168;
razn_w_mem[12335] = 168;
razn_w_mem[12336] = 168;
razn_w_mem[12337] = 168;
razn_w_mem[12338] = 168;
razn_w_mem[12339] = 168;
razn_w_mem[12340] = 168;
razn_w_mem[12341] = 168;
razn_w_mem[12342] = 168;
razn_w_mem[12343] = 168;
razn_w_mem[12344] = 168;
razn_w_mem[12345] = 168;
razn_w_mem[12346] = 168;
razn_w_mem[12347] = 168;
razn_w_mem[12348] = 168;
razn_w_mem[12349] = 168;
razn_w_mem[12350] = 168;
razn_w_mem[12351] = 168;
razn_w_mem[12352] = 168;
razn_w_mem[12353] = 168;
razn_w_mem[12354] = 168;
razn_w_mem[12355] = 168;
razn_w_mem[12356] = 168;
razn_w_mem[12357] = 168;
razn_w_mem[12358] = 168;
razn_w_mem[12359] = 168;
razn_w_mem[12360] = 168;
razn_w_mem[12361] = 168;
razn_w_mem[12362] = 168;
razn_w_mem[12363] = 168;
razn_w_mem[12364] = 168;
razn_w_mem[12365] = 168;
razn_w_mem[12366] = 168;
razn_w_mem[12367] = 168;
razn_w_mem[12368] = 168;
razn_w_mem[12369] = 168;
razn_w_mem[12370] = 168;
razn_w_mem[12371] = 168;
razn_w_mem[12372] = 168;
razn_w_mem[12373] = 168;
razn_w_mem[12374] = 168;
razn_w_mem[12375] = 168;
razn_w_mem[12376] = 168;
razn_w_mem[12377] = 168;
razn_w_mem[12378] = 168;
razn_w_mem[12379] = 168;
razn_w_mem[12380] = 168;
razn_w_mem[12381] = 168;
razn_w_mem[12382] = 168;
razn_w_mem[12383] = 168;
razn_w_mem[12384] = 168;
razn_w_mem[12385] = 168;
razn_w_mem[12386] = 168;
razn_w_mem[12387] = 168;
razn_w_mem[12388] = 168;
razn_w_mem[12389] = 168;
razn_w_mem[12390] = 168;
razn_w_mem[12391] = 168;
razn_w_mem[12392] = 168;
razn_w_mem[12393] = 168;
razn_w_mem[12394] = 168;
razn_w_mem[12395] = 168;
razn_w_mem[12396] = 168;
razn_w_mem[12397] = 168;
razn_w_mem[12398] = 168;
razn_w_mem[12399] = 168;
razn_w_mem[12400] = 168;
razn_w_mem[12401] = 168;
razn_w_mem[12402] = 168;
razn_w_mem[12403] = 168;
razn_w_mem[12404] = 168;
razn_w_mem[12405] = 168;
razn_w_mem[12406] = 168;
razn_w_mem[12407] = 168;
razn_w_mem[12408] = 168;
razn_w_mem[12409] = 168;
razn_w_mem[12410] = 168;
razn_w_mem[12411] = 168;
razn_w_mem[12412] = 168;
razn_w_mem[12413] = 168;
razn_w_mem[12414] = 168;
razn_w_mem[12415] = 168;
razn_w_mem[12416] = 138;
razn_w_mem[12417] = 138;
razn_w_mem[12418] = 138;
razn_w_mem[12419] = 138;
razn_w_mem[12420] = 138;
razn_w_mem[12421] = 138;
razn_w_mem[12422] = 138;
razn_w_mem[12423] = 138;
razn_w_mem[12424] = 138;
razn_w_mem[12425] = 138;
razn_w_mem[12426] = 138;
razn_w_mem[12427] = 138;
razn_w_mem[12428] = 138;
razn_w_mem[12429] = 138;
razn_w_mem[12430] = 138;
razn_w_mem[12431] = 138;
razn_w_mem[12432] = 138;
razn_w_mem[12433] = 138;
razn_w_mem[12434] = 138;
razn_w_mem[12435] = 138;
razn_w_mem[12436] = 138;
razn_w_mem[12437] = 138;
razn_w_mem[12438] = 138;
razn_w_mem[12439] = 138;
razn_w_mem[12440] = 138;
razn_w_mem[12441] = 138;
razn_w_mem[12442] = 138;
razn_w_mem[12443] = 138;
razn_w_mem[12444] = 138;
razn_w_mem[12445] = 138;
razn_w_mem[12446] = 138;
razn_w_mem[12447] = 138;
razn_w_mem[12448] = 138;
razn_w_mem[12449] = 138;
razn_w_mem[12450] = 138;
razn_w_mem[12451] = 138;
razn_w_mem[12452] = 138;
razn_w_mem[12453] = 138;
razn_w_mem[12454] = 138;
razn_w_mem[12455] = 138;
razn_w_mem[12456] = 138;
razn_w_mem[12457] = 138;
razn_w_mem[12458] = 138;
razn_w_mem[12459] = 138;
razn_w_mem[12460] = 138;
razn_w_mem[12461] = 138;
razn_w_mem[12462] = 138;
razn_w_mem[12463] = 138;
razn_w_mem[12464] = 138;
razn_w_mem[12465] = 138;
razn_w_mem[12466] = 138;
razn_w_mem[12467] = 138;
razn_w_mem[12468] = 138;
razn_w_mem[12469] = 138;
razn_w_mem[12470] = 138;
razn_w_mem[12471] = 138;
razn_w_mem[12472] = 138;
razn_w_mem[12473] = 138;
razn_w_mem[12474] = 138;
razn_w_mem[12475] = 138;
razn_w_mem[12476] = 138;
razn_w_mem[12477] = 138;
razn_w_mem[12478] = 138;
razn_w_mem[12479] = 138;
razn_w_mem[12480] = 138;
razn_w_mem[12481] = 138;
razn_w_mem[12482] = 138;
razn_w_mem[12483] = 138;
razn_w_mem[12484] = 138;
razn_w_mem[12485] = 138;
razn_w_mem[12486] = 138;
razn_w_mem[12487] = 138;
razn_w_mem[12488] = 138;
razn_w_mem[12489] = 138;
razn_w_mem[12490] = 138;
razn_w_mem[12491] = 138;
razn_w_mem[12492] = 138;
razn_w_mem[12493] = 138;
razn_w_mem[12494] = 138;
razn_w_mem[12495] = 138;
razn_w_mem[12496] = 138;
razn_w_mem[12497] = 138;
razn_w_mem[12498] = 138;
razn_w_mem[12499] = 138;
razn_w_mem[12500] = 138;
razn_w_mem[12501] = 138;
razn_w_mem[12502] = 138;
razn_w_mem[12503] = 138;
razn_w_mem[12504] = 138;
razn_w_mem[12505] = 138;
razn_w_mem[12506] = 138;
razn_w_mem[12507] = 138;
razn_w_mem[12508] = 138;
razn_w_mem[12509] = 138;
razn_w_mem[12510] = 138;
razn_w_mem[12511] = 138;
razn_w_mem[12512] = 138;
razn_w_mem[12513] = 138;
razn_w_mem[12514] = 138;
razn_w_mem[12515] = 138;
razn_w_mem[12516] = 138;
razn_w_mem[12517] = 138;
razn_w_mem[12518] = 138;
razn_w_mem[12519] = 138;
razn_w_mem[12520] = 138;
razn_w_mem[12521] = 138;
razn_w_mem[12522] = 138;
razn_w_mem[12523] = 138;
razn_w_mem[12524] = 138;
razn_w_mem[12525] = 138;
razn_w_mem[12526] = 138;
razn_w_mem[12527] = 138;
razn_w_mem[12528] = 138;
razn_w_mem[12529] = 138;
razn_w_mem[12530] = 138;
razn_w_mem[12531] = 138;
razn_w_mem[12532] = 138;
razn_w_mem[12533] = 138;
razn_w_mem[12534] = 138;
razn_w_mem[12535] = 138;
razn_w_mem[12536] = 138;
razn_w_mem[12537] = 138;
razn_w_mem[12538] = 138;
razn_w_mem[12539] = 138;
razn_w_mem[12540] = 138;
razn_w_mem[12541] = 138;
razn_w_mem[12542] = 138;
razn_w_mem[12543] = 138;
razn_w_mem[12544] = 108;
razn_w_mem[12545] = 108;
razn_w_mem[12546] = 108;
razn_w_mem[12547] = 108;
razn_w_mem[12548] = 108;
razn_w_mem[12549] = 108;
razn_w_mem[12550] = 108;
razn_w_mem[12551] = 108;
razn_w_mem[12552] = 108;
razn_w_mem[12553] = 108;
razn_w_mem[12554] = 108;
razn_w_mem[12555] = 108;
razn_w_mem[12556] = 108;
razn_w_mem[12557] = 108;
razn_w_mem[12558] = 108;
razn_w_mem[12559] = 108;
razn_w_mem[12560] = 108;
razn_w_mem[12561] = 108;
razn_w_mem[12562] = 108;
razn_w_mem[12563] = 108;
razn_w_mem[12564] = 108;
razn_w_mem[12565] = 108;
razn_w_mem[12566] = 108;
razn_w_mem[12567] = 108;
razn_w_mem[12568] = 108;
razn_w_mem[12569] = 108;
razn_w_mem[12570] = 108;
razn_w_mem[12571] = 108;
razn_w_mem[12572] = 108;
razn_w_mem[12573] = 108;
razn_w_mem[12574] = 108;
razn_w_mem[12575] = 108;
razn_w_mem[12576] = 108;
razn_w_mem[12577] = 108;
razn_w_mem[12578] = 108;
razn_w_mem[12579] = 108;
razn_w_mem[12580] = 108;
razn_w_mem[12581] = 108;
razn_w_mem[12582] = 108;
razn_w_mem[12583] = 108;
razn_w_mem[12584] = 108;
razn_w_mem[12585] = 108;
razn_w_mem[12586] = 108;
razn_w_mem[12587] = 108;
razn_w_mem[12588] = 108;
razn_w_mem[12589] = 108;
razn_w_mem[12590] = 108;
razn_w_mem[12591] = 108;
razn_w_mem[12592] = 108;
razn_w_mem[12593] = 108;
razn_w_mem[12594] = 108;
razn_w_mem[12595] = 108;
razn_w_mem[12596] = 108;
razn_w_mem[12597] = 108;
razn_w_mem[12598] = 108;
razn_w_mem[12599] = 108;
razn_w_mem[12600] = 108;
razn_w_mem[12601] = 108;
razn_w_mem[12602] = 108;
razn_w_mem[12603] = 108;
razn_w_mem[12604] = 108;
razn_w_mem[12605] = 108;
razn_w_mem[12606] = 108;
razn_w_mem[12607] = 108;
razn_w_mem[12608] = 108;
razn_w_mem[12609] = 108;
razn_w_mem[12610] = 108;
razn_w_mem[12611] = 108;
razn_w_mem[12612] = 108;
razn_w_mem[12613] = 108;
razn_w_mem[12614] = 108;
razn_w_mem[12615] = 108;
razn_w_mem[12616] = 108;
razn_w_mem[12617] = 108;
razn_w_mem[12618] = 108;
razn_w_mem[12619] = 108;
razn_w_mem[12620] = 108;
razn_w_mem[12621] = 108;
razn_w_mem[12622] = 108;
razn_w_mem[12623] = 108;
razn_w_mem[12624] = 108;
razn_w_mem[12625] = 108;
razn_w_mem[12626] = 108;
razn_w_mem[12627] = 108;
razn_w_mem[12628] = 108;
razn_w_mem[12629] = 108;
razn_w_mem[12630] = 108;
razn_w_mem[12631] = 108;
razn_w_mem[12632] = 108;
razn_w_mem[12633] = 108;
razn_w_mem[12634] = 108;
razn_w_mem[12635] = 108;
razn_w_mem[12636] = 108;
razn_w_mem[12637] = 108;
razn_w_mem[12638] = 108;
razn_w_mem[12639] = 108;
razn_w_mem[12640] = 108;
razn_w_mem[12641] = 108;
razn_w_mem[12642] = 108;
razn_w_mem[12643] = 108;
razn_w_mem[12644] = 108;
razn_w_mem[12645] = 108;
razn_w_mem[12646] = 108;
razn_w_mem[12647] = 108;
razn_w_mem[12648] = 108;
razn_w_mem[12649] = 108;
razn_w_mem[12650] = 108;
razn_w_mem[12651] = 108;
razn_w_mem[12652] = 108;
razn_w_mem[12653] = 108;
razn_w_mem[12654] = 108;
razn_w_mem[12655] = 108;
razn_w_mem[12656] = 108;
razn_w_mem[12657] = 108;
razn_w_mem[12658] = 108;
razn_w_mem[12659] = 108;
razn_w_mem[12660] = 108;
razn_w_mem[12661] = 108;
razn_w_mem[12662] = 108;
razn_w_mem[12663] = 108;
razn_w_mem[12664] = 108;
razn_w_mem[12665] = 108;
razn_w_mem[12666] = 108;
razn_w_mem[12667] = 108;
razn_w_mem[12668] = 108;
razn_w_mem[12669] = 108;
razn_w_mem[12670] = 108;
razn_w_mem[12671] = 108;
razn_w_mem[12672] = 78;
razn_w_mem[12673] = 78;
razn_w_mem[12674] = 78;
razn_w_mem[12675] = 78;
razn_w_mem[12676] = 78;
razn_w_mem[12677] = 78;
razn_w_mem[12678] = 78;
razn_w_mem[12679] = 78;
razn_w_mem[12680] = 78;
razn_w_mem[12681] = 78;
razn_w_mem[12682] = 78;
razn_w_mem[12683] = 78;
razn_w_mem[12684] = 78;
razn_w_mem[12685] = 78;
razn_w_mem[12686] = 78;
razn_w_mem[12687] = 78;
razn_w_mem[12688] = 78;
razn_w_mem[12689] = 78;
razn_w_mem[12690] = 78;
razn_w_mem[12691] = 78;
razn_w_mem[12692] = 78;
razn_w_mem[12693] = 78;
razn_w_mem[12694] = 78;
razn_w_mem[12695] = 78;
razn_w_mem[12696] = 78;
razn_w_mem[12697] = 78;
razn_w_mem[12698] = 78;
razn_w_mem[12699] = 78;
razn_w_mem[12700] = 78;
razn_w_mem[12701] = 78;
razn_w_mem[12702] = 78;
razn_w_mem[12703] = 78;
razn_w_mem[12704] = 78;
razn_w_mem[12705] = 78;
razn_w_mem[12706] = 78;
razn_w_mem[12707] = 78;
razn_w_mem[12708] = 78;
razn_w_mem[12709] = 78;
razn_w_mem[12710] = 78;
razn_w_mem[12711] = 78;
razn_w_mem[12712] = 78;
razn_w_mem[12713] = 78;
razn_w_mem[12714] = 78;
razn_w_mem[12715] = 78;
razn_w_mem[12716] = 78;
razn_w_mem[12717] = 78;
razn_w_mem[12718] = 78;
razn_w_mem[12719] = 78;
razn_w_mem[12720] = 78;
razn_w_mem[12721] = 78;
razn_w_mem[12722] = 78;
razn_w_mem[12723] = 78;
razn_w_mem[12724] = 78;
razn_w_mem[12725] = 78;
razn_w_mem[12726] = 78;
razn_w_mem[12727] = 78;
razn_w_mem[12728] = 78;
razn_w_mem[12729] = 78;
razn_w_mem[12730] = 78;
razn_w_mem[12731] = 78;
razn_w_mem[12732] = 78;
razn_w_mem[12733] = 78;
razn_w_mem[12734] = 78;
razn_w_mem[12735] = 78;
razn_w_mem[12736] = 78;
razn_w_mem[12737] = 78;
razn_w_mem[12738] = 78;
razn_w_mem[12739] = 78;
razn_w_mem[12740] = 78;
razn_w_mem[12741] = 78;
razn_w_mem[12742] = 78;
razn_w_mem[12743] = 78;
razn_w_mem[12744] = 78;
razn_w_mem[12745] = 78;
razn_w_mem[12746] = 78;
razn_w_mem[12747] = 78;
razn_w_mem[12748] = 78;
razn_w_mem[12749] = 78;
razn_w_mem[12750] = 78;
razn_w_mem[12751] = 78;
razn_w_mem[12752] = 78;
razn_w_mem[12753] = 78;
razn_w_mem[12754] = 78;
razn_w_mem[12755] = 78;
razn_w_mem[12756] = 78;
razn_w_mem[12757] = 78;
razn_w_mem[12758] = 78;
razn_w_mem[12759] = 78;
razn_w_mem[12760] = 78;
razn_w_mem[12761] = 78;
razn_w_mem[12762] = 78;
razn_w_mem[12763] = 78;
razn_w_mem[12764] = 78;
razn_w_mem[12765] = 78;
razn_w_mem[12766] = 78;
razn_w_mem[12767] = 78;
razn_w_mem[12768] = 78;
razn_w_mem[12769] = 78;
razn_w_mem[12770] = 78;
razn_w_mem[12771] = 78;
razn_w_mem[12772] = 78;
razn_w_mem[12773] = 78;
razn_w_mem[12774] = 78;
razn_w_mem[12775] = 78;
razn_w_mem[12776] = 78;
razn_w_mem[12777] = 78;
razn_w_mem[12778] = 78;
razn_w_mem[12779] = 78;
razn_w_mem[12780] = 78;
razn_w_mem[12781] = 78;
razn_w_mem[12782] = 78;
razn_w_mem[12783] = 78;
razn_w_mem[12784] = 78;
razn_w_mem[12785] = 78;
razn_w_mem[12786] = 78;
razn_w_mem[12787] = 78;
razn_w_mem[12788] = 78;
razn_w_mem[12789] = 78;
razn_w_mem[12790] = 78;
razn_w_mem[12791] = 78;
razn_w_mem[12792] = 78;
razn_w_mem[12793] = 78;
razn_w_mem[12794] = 78;
razn_w_mem[12795] = 78;
razn_w_mem[12796] = 78;
razn_w_mem[12797] = 78;
razn_w_mem[12798] = 78;
razn_w_mem[12799] = 78;
razn_w_mem[12800] = 48;
razn_w_mem[12801] = 48;
razn_w_mem[12802] = 48;
razn_w_mem[12803] = 48;
razn_w_mem[12804] = 48;
razn_w_mem[12805] = 48;
razn_w_mem[12806] = 48;
razn_w_mem[12807] = 48;
razn_w_mem[12808] = 48;
razn_w_mem[12809] = 48;
razn_w_mem[12810] = 48;
razn_w_mem[12811] = 48;
razn_w_mem[12812] = 48;
razn_w_mem[12813] = 48;
razn_w_mem[12814] = 48;
razn_w_mem[12815] = 48;
razn_w_mem[12816] = 48;
razn_w_mem[12817] = 48;
razn_w_mem[12818] = 48;
razn_w_mem[12819] = 48;
razn_w_mem[12820] = 48;
razn_w_mem[12821] = 48;
razn_w_mem[12822] = 48;
razn_w_mem[12823] = 48;
razn_w_mem[12824] = 48;
razn_w_mem[12825] = 48;
razn_w_mem[12826] = 48;
razn_w_mem[12827] = 48;
razn_w_mem[12828] = 48;
razn_w_mem[12829] = 48;
razn_w_mem[12830] = 48;
razn_w_mem[12831] = 48;
razn_w_mem[12832] = 48;
razn_w_mem[12833] = 48;
razn_w_mem[12834] = 48;
razn_w_mem[12835] = 48;
razn_w_mem[12836] = 48;
razn_w_mem[12837] = 48;
razn_w_mem[12838] = 48;
razn_w_mem[12839] = 48;
razn_w_mem[12840] = 48;
razn_w_mem[12841] = 48;
razn_w_mem[12842] = 48;
razn_w_mem[12843] = 48;
razn_w_mem[12844] = 48;
razn_w_mem[12845] = 48;
razn_w_mem[12846] = 48;
razn_w_mem[12847] = 48;
razn_w_mem[12848] = 48;
razn_w_mem[12849] = 48;
razn_w_mem[12850] = 48;
razn_w_mem[12851] = 48;
razn_w_mem[12852] = 48;
razn_w_mem[12853] = 48;
razn_w_mem[12854] = 48;
razn_w_mem[12855] = 48;
razn_w_mem[12856] = 48;
razn_w_mem[12857] = 48;
razn_w_mem[12858] = 48;
razn_w_mem[12859] = 48;
razn_w_mem[12860] = 48;
razn_w_mem[12861] = 48;
razn_w_mem[12862] = 48;
razn_w_mem[12863] = 48;
razn_w_mem[12864] = 48;
razn_w_mem[12865] = 48;
razn_w_mem[12866] = 48;
razn_w_mem[12867] = 48;
razn_w_mem[12868] = 48;
razn_w_mem[12869] = 48;
razn_w_mem[12870] = 48;
razn_w_mem[12871] = 48;
razn_w_mem[12872] = 48;
razn_w_mem[12873] = 48;
razn_w_mem[12874] = 48;
razn_w_mem[12875] = 48;
razn_w_mem[12876] = 48;
razn_w_mem[12877] = 48;
razn_w_mem[12878] = 48;
razn_w_mem[12879] = 48;
razn_w_mem[12880] = 48;
razn_w_mem[12881] = 48;
razn_w_mem[12882] = 48;
razn_w_mem[12883] = 48;
razn_w_mem[12884] = 48;
razn_w_mem[12885] = 48;
razn_w_mem[12886] = 48;
razn_w_mem[12887] = 48;
razn_w_mem[12888] = 48;
razn_w_mem[12889] = 48;
razn_w_mem[12890] = 48;
razn_w_mem[12891] = 48;
razn_w_mem[12892] = 48;
razn_w_mem[12893] = 48;
razn_w_mem[12894] = 48;
razn_w_mem[12895] = 48;
razn_w_mem[12896] = 48;
razn_w_mem[12897] = 48;
razn_w_mem[12898] = 48;
razn_w_mem[12899] = 48;
razn_w_mem[12900] = 48;
razn_w_mem[12901] = 48;
razn_w_mem[12902] = 48;
razn_w_mem[12903] = 48;
razn_w_mem[12904] = 48;
razn_w_mem[12905] = 48;
razn_w_mem[12906] = 48;
razn_w_mem[12907] = 48;
razn_w_mem[12908] = 48;
razn_w_mem[12909] = 48;
razn_w_mem[12910] = 48;
razn_w_mem[12911] = 48;
razn_w_mem[12912] = 48;
razn_w_mem[12913] = 48;
razn_w_mem[12914] = 48;
razn_w_mem[12915] = 48;
razn_w_mem[12916] = 48;
razn_w_mem[12917] = 48;
razn_w_mem[12918] = 48;
razn_w_mem[12919] = 48;
razn_w_mem[12920] = 48;
razn_w_mem[12921] = 48;
razn_w_mem[12922] = 48;
razn_w_mem[12923] = 48;
razn_w_mem[12924] = 48;
razn_w_mem[12925] = 48;
razn_w_mem[12926] = 48;
razn_w_mem[12927] = 48;
razn_w_mem[12928] = 18;
razn_w_mem[12929] = 18;
razn_w_mem[12930] = 18;
razn_w_mem[12931] = 18;
razn_w_mem[12932] = 18;
razn_w_mem[12933] = 18;
razn_w_mem[12934] = 18;
razn_w_mem[12935] = 18;
razn_w_mem[12936] = 18;
razn_w_mem[12937] = 18;
razn_w_mem[12938] = 18;
razn_w_mem[12939] = 18;
razn_w_mem[12940] = 18;
razn_w_mem[12941] = 18;
razn_w_mem[12942] = 18;
razn_w_mem[12943] = 18;
razn_w_mem[12944] = 18;
razn_w_mem[12945] = 18;
razn_w_mem[12946] = 18;
razn_w_mem[12947] = 18;
razn_w_mem[12948] = 18;
razn_w_mem[12949] = 18;
razn_w_mem[12950] = 18;
razn_w_mem[12951] = 18;
razn_w_mem[12952] = 18;
razn_w_mem[12953] = 18;
razn_w_mem[12954] = 18;
razn_w_mem[12955] = 18;
razn_w_mem[12956] = 18;
razn_w_mem[12957] = 18;
razn_w_mem[12958] = 18;
razn_w_mem[12959] = 18;
razn_w_mem[12960] = 18;
razn_w_mem[12961] = 18;
razn_w_mem[12962] = 18;
razn_w_mem[12963] = 18;
razn_w_mem[12964] = 18;
razn_w_mem[12965] = 18;
razn_w_mem[12966] = 18;
razn_w_mem[12967] = 18;
razn_w_mem[12968] = 18;
razn_w_mem[12969] = 18;
razn_w_mem[12970] = 18;
razn_w_mem[12971] = 18;
razn_w_mem[12972] = 18;
razn_w_mem[12973] = 18;
razn_w_mem[12974] = 18;
razn_w_mem[12975] = 18;
razn_w_mem[12976] = 18;
razn_w_mem[12977] = 18;
razn_w_mem[12978] = 18;
razn_w_mem[12979] = 18;
razn_w_mem[12980] = 18;
razn_w_mem[12981] = 18;
razn_w_mem[12982] = 18;
razn_w_mem[12983] = 18;
razn_w_mem[12984] = 18;
razn_w_mem[12985] = 18;
razn_w_mem[12986] = 18;
razn_w_mem[12987] = 18;
razn_w_mem[12988] = 18;
razn_w_mem[12989] = 18;
razn_w_mem[12990] = 18;
razn_w_mem[12991] = 18;
razn_w_mem[12992] = 18;
razn_w_mem[12993] = 18;
razn_w_mem[12994] = 18;
razn_w_mem[12995] = 18;
razn_w_mem[12996] = 18;
razn_w_mem[12997] = 18;
razn_w_mem[12998] = 18;
razn_w_mem[12999] = 18;
razn_w_mem[13000] = 18;
razn_w_mem[13001] = 18;
razn_w_mem[13002] = 18;
razn_w_mem[13003] = 18;
razn_w_mem[13004] = 18;
razn_w_mem[13005] = 18;
razn_w_mem[13006] = 18;
razn_w_mem[13007] = 18;
razn_w_mem[13008] = 18;
razn_w_mem[13009] = 18;
razn_w_mem[13010] = 18;
razn_w_mem[13011] = 18;
razn_w_mem[13012] = 18;
razn_w_mem[13013] = 18;
razn_w_mem[13014] = 18;
razn_w_mem[13015] = 18;
razn_w_mem[13016] = 18;
razn_w_mem[13017] = 18;
razn_w_mem[13018] = 18;
razn_w_mem[13019] = 18;
razn_w_mem[13020] = 18;
razn_w_mem[13021] = 18;
razn_w_mem[13022] = 18;
razn_w_mem[13023] = 18;
razn_w_mem[13024] = 18;
razn_w_mem[13025] = 18;
razn_w_mem[13026] = 18;
razn_w_mem[13027] = 18;
razn_w_mem[13028] = 18;
razn_w_mem[13029] = 18;
razn_w_mem[13030] = 18;
razn_w_mem[13031] = 18;
razn_w_mem[13032] = 18;
razn_w_mem[13033] = 18;
razn_w_mem[13034] = 18;
razn_w_mem[13035] = 18;
razn_w_mem[13036] = 18;
razn_w_mem[13037] = 18;
razn_w_mem[13038] = 18;
razn_w_mem[13039] = 18;
razn_w_mem[13040] = 18;
razn_w_mem[13041] = 18;
razn_w_mem[13042] = 18;
razn_w_mem[13043] = 18;
razn_w_mem[13044] = 18;
razn_w_mem[13045] = 18;
razn_w_mem[13046] = 18;
razn_w_mem[13047] = 18;
razn_w_mem[13048] = 18;
razn_w_mem[13049] = 18;
razn_w_mem[13050] = 18;
razn_w_mem[13051] = 18;
razn_w_mem[13052] = 18;
razn_w_mem[13053] = 18;
razn_w_mem[13054] = 18;
razn_w_mem[13055] = 18;
razn_w_mem[13056] = 242;
razn_w_mem[13057] = 242;
razn_w_mem[13058] = 242;
razn_w_mem[13059] = 242;
razn_w_mem[13060] = 242;
razn_w_mem[13061] = 242;
razn_w_mem[13062] = 242;
razn_w_mem[13063] = 242;
razn_w_mem[13064] = 242;
razn_w_mem[13065] = 242;
razn_w_mem[13066] = 242;
razn_w_mem[13067] = 242;
razn_w_mem[13068] = 242;
razn_w_mem[13069] = 242;
razn_w_mem[13070] = 242;
razn_w_mem[13071] = 242;
razn_w_mem[13072] = 242;
razn_w_mem[13073] = 242;
razn_w_mem[13074] = 242;
razn_w_mem[13075] = 242;
razn_w_mem[13076] = 242;
razn_w_mem[13077] = 242;
razn_w_mem[13078] = 242;
razn_w_mem[13079] = 242;
razn_w_mem[13080] = 242;
razn_w_mem[13081] = 242;
razn_w_mem[13082] = 242;
razn_w_mem[13083] = 242;
razn_w_mem[13084] = 242;
razn_w_mem[13085] = 242;
razn_w_mem[13086] = 242;
razn_w_mem[13087] = 242;
razn_w_mem[13088] = 242;
razn_w_mem[13089] = 242;
razn_w_mem[13090] = 242;
razn_w_mem[13091] = 242;
razn_w_mem[13092] = 242;
razn_w_mem[13093] = 242;
razn_w_mem[13094] = 242;
razn_w_mem[13095] = 242;
razn_w_mem[13096] = 242;
razn_w_mem[13097] = 242;
razn_w_mem[13098] = 242;
razn_w_mem[13099] = 242;
razn_w_mem[13100] = 242;
razn_w_mem[13101] = 242;
razn_w_mem[13102] = 242;
razn_w_mem[13103] = 242;
razn_w_mem[13104] = 242;
razn_w_mem[13105] = 242;
razn_w_mem[13106] = 242;
razn_w_mem[13107] = 242;
razn_w_mem[13108] = 242;
razn_w_mem[13109] = 242;
razn_w_mem[13110] = 242;
razn_w_mem[13111] = 242;
razn_w_mem[13112] = 242;
razn_w_mem[13113] = 242;
razn_w_mem[13114] = 242;
razn_w_mem[13115] = 242;
razn_w_mem[13116] = 242;
razn_w_mem[13117] = 242;
razn_w_mem[13118] = 242;
razn_w_mem[13119] = 242;
razn_w_mem[13120] = 242;
razn_w_mem[13121] = 242;
razn_w_mem[13122] = 242;
razn_w_mem[13123] = 242;
razn_w_mem[13124] = 242;
razn_w_mem[13125] = 242;
razn_w_mem[13126] = 242;
razn_w_mem[13127] = 242;
razn_w_mem[13128] = 242;
razn_w_mem[13129] = 242;
razn_w_mem[13130] = 242;
razn_w_mem[13131] = 242;
razn_w_mem[13132] = 242;
razn_w_mem[13133] = 242;
razn_w_mem[13134] = 242;
razn_w_mem[13135] = 242;
razn_w_mem[13136] = 242;
razn_w_mem[13137] = 242;
razn_w_mem[13138] = 242;
razn_w_mem[13139] = 242;
razn_w_mem[13140] = 242;
razn_w_mem[13141] = 242;
razn_w_mem[13142] = 242;
razn_w_mem[13143] = 242;
razn_w_mem[13144] = 242;
razn_w_mem[13145] = 242;
razn_w_mem[13146] = 242;
razn_w_mem[13147] = 242;
razn_w_mem[13148] = 242;
razn_w_mem[13149] = 242;
razn_w_mem[13150] = 242;
razn_w_mem[13151] = 242;
razn_w_mem[13152] = 242;
razn_w_mem[13153] = 242;
razn_w_mem[13154] = 242;
razn_w_mem[13155] = 242;
razn_w_mem[13156] = 242;
razn_w_mem[13157] = 242;
razn_w_mem[13158] = 242;
razn_w_mem[13159] = 242;
razn_w_mem[13160] = 242;
razn_w_mem[13161] = 242;
razn_w_mem[13162] = 242;
razn_w_mem[13163] = 242;
razn_w_mem[13164] = 242;
razn_w_mem[13165] = 242;
razn_w_mem[13166] = 242;
razn_w_mem[13167] = 242;
razn_w_mem[13168] = 242;
razn_w_mem[13169] = 242;
razn_w_mem[13170] = 242;
razn_w_mem[13171] = 242;
razn_w_mem[13172] = 242;
razn_w_mem[13173] = 242;
razn_w_mem[13174] = 242;
razn_w_mem[13175] = 242;
razn_w_mem[13176] = 242;
razn_w_mem[13177] = 242;
razn_w_mem[13178] = 242;
razn_w_mem[13179] = 242;
razn_w_mem[13180] = 242;
razn_w_mem[13181] = 242;
razn_w_mem[13182] = 242;
razn_w_mem[13183] = 242;
razn_w_mem[13184] = 212;
razn_w_mem[13185] = 212;
razn_w_mem[13186] = 212;
razn_w_mem[13187] = 212;
razn_w_mem[13188] = 212;
razn_w_mem[13189] = 212;
razn_w_mem[13190] = 212;
razn_w_mem[13191] = 212;
razn_w_mem[13192] = 212;
razn_w_mem[13193] = 212;
razn_w_mem[13194] = 212;
razn_w_mem[13195] = 212;
razn_w_mem[13196] = 212;
razn_w_mem[13197] = 212;
razn_w_mem[13198] = 212;
razn_w_mem[13199] = 212;
razn_w_mem[13200] = 212;
razn_w_mem[13201] = 212;
razn_w_mem[13202] = 212;
razn_w_mem[13203] = 212;
razn_w_mem[13204] = 212;
razn_w_mem[13205] = 212;
razn_w_mem[13206] = 212;
razn_w_mem[13207] = 212;
razn_w_mem[13208] = 212;
razn_w_mem[13209] = 212;
razn_w_mem[13210] = 212;
razn_w_mem[13211] = 212;
razn_w_mem[13212] = 212;
razn_w_mem[13213] = 212;
razn_w_mem[13214] = 212;
razn_w_mem[13215] = 212;
razn_w_mem[13216] = 212;
razn_w_mem[13217] = 212;
razn_w_mem[13218] = 212;
razn_w_mem[13219] = 212;
razn_w_mem[13220] = 212;
razn_w_mem[13221] = 212;
razn_w_mem[13222] = 212;
razn_w_mem[13223] = 212;
razn_w_mem[13224] = 212;
razn_w_mem[13225] = 212;
razn_w_mem[13226] = 212;
razn_w_mem[13227] = 212;
razn_w_mem[13228] = 212;
razn_w_mem[13229] = 212;
razn_w_mem[13230] = 212;
razn_w_mem[13231] = 212;
razn_w_mem[13232] = 212;
razn_w_mem[13233] = 212;
razn_w_mem[13234] = 212;
razn_w_mem[13235] = 212;
razn_w_mem[13236] = 212;
razn_w_mem[13237] = 212;
razn_w_mem[13238] = 212;
razn_w_mem[13239] = 212;
razn_w_mem[13240] = 212;
razn_w_mem[13241] = 212;
razn_w_mem[13242] = 212;
razn_w_mem[13243] = 212;
razn_w_mem[13244] = 212;
razn_w_mem[13245] = 212;
razn_w_mem[13246] = 212;
razn_w_mem[13247] = 212;
razn_w_mem[13248] = 212;
razn_w_mem[13249] = 212;
razn_w_mem[13250] = 212;
razn_w_mem[13251] = 212;
razn_w_mem[13252] = 212;
razn_w_mem[13253] = 212;
razn_w_mem[13254] = 212;
razn_w_mem[13255] = 212;
razn_w_mem[13256] = 212;
razn_w_mem[13257] = 212;
razn_w_mem[13258] = 212;
razn_w_mem[13259] = 212;
razn_w_mem[13260] = 212;
razn_w_mem[13261] = 212;
razn_w_mem[13262] = 212;
razn_w_mem[13263] = 212;
razn_w_mem[13264] = 212;
razn_w_mem[13265] = 212;
razn_w_mem[13266] = 212;
razn_w_mem[13267] = 212;
razn_w_mem[13268] = 212;
razn_w_mem[13269] = 212;
razn_w_mem[13270] = 212;
razn_w_mem[13271] = 212;
razn_w_mem[13272] = 212;
razn_w_mem[13273] = 212;
razn_w_mem[13274] = 212;
razn_w_mem[13275] = 212;
razn_w_mem[13276] = 212;
razn_w_mem[13277] = 212;
razn_w_mem[13278] = 212;
razn_w_mem[13279] = 212;
razn_w_mem[13280] = 212;
razn_w_mem[13281] = 212;
razn_w_mem[13282] = 212;
razn_w_mem[13283] = 212;
razn_w_mem[13284] = 212;
razn_w_mem[13285] = 212;
razn_w_mem[13286] = 212;
razn_w_mem[13287] = 212;
razn_w_mem[13288] = 212;
razn_w_mem[13289] = 212;
razn_w_mem[13290] = 212;
razn_w_mem[13291] = 212;
razn_w_mem[13292] = 212;
razn_w_mem[13293] = 212;
razn_w_mem[13294] = 212;
razn_w_mem[13295] = 212;
razn_w_mem[13296] = 212;
razn_w_mem[13297] = 212;
razn_w_mem[13298] = 212;
razn_w_mem[13299] = 212;
razn_w_mem[13300] = 212;
razn_w_mem[13301] = 212;
razn_w_mem[13302] = 212;
razn_w_mem[13303] = 212;
razn_w_mem[13304] = 212;
razn_w_mem[13305] = 212;
razn_w_mem[13306] = 212;
razn_w_mem[13307] = 212;
razn_w_mem[13308] = 212;
razn_w_mem[13309] = 212;
razn_w_mem[13310] = 212;
razn_w_mem[13311] = 212;
razn_w_mem[13312] = 182;
razn_w_mem[13313] = 182;
razn_w_mem[13314] = 182;
razn_w_mem[13315] = 182;
razn_w_mem[13316] = 182;
razn_w_mem[13317] = 182;
razn_w_mem[13318] = 182;
razn_w_mem[13319] = 182;
razn_w_mem[13320] = 182;
razn_w_mem[13321] = 182;
razn_w_mem[13322] = 182;
razn_w_mem[13323] = 182;
razn_w_mem[13324] = 182;
razn_w_mem[13325] = 182;
razn_w_mem[13326] = 182;
razn_w_mem[13327] = 182;
razn_w_mem[13328] = 182;
razn_w_mem[13329] = 182;
razn_w_mem[13330] = 182;
razn_w_mem[13331] = 182;
razn_w_mem[13332] = 182;
razn_w_mem[13333] = 182;
razn_w_mem[13334] = 182;
razn_w_mem[13335] = 182;
razn_w_mem[13336] = 182;
razn_w_mem[13337] = 182;
razn_w_mem[13338] = 182;
razn_w_mem[13339] = 182;
razn_w_mem[13340] = 182;
razn_w_mem[13341] = 182;
razn_w_mem[13342] = 182;
razn_w_mem[13343] = 182;
razn_w_mem[13344] = 182;
razn_w_mem[13345] = 182;
razn_w_mem[13346] = 182;
razn_w_mem[13347] = 182;
razn_w_mem[13348] = 182;
razn_w_mem[13349] = 182;
razn_w_mem[13350] = 182;
razn_w_mem[13351] = 182;
razn_w_mem[13352] = 182;
razn_w_mem[13353] = 182;
razn_w_mem[13354] = 182;
razn_w_mem[13355] = 182;
razn_w_mem[13356] = 182;
razn_w_mem[13357] = 182;
razn_w_mem[13358] = 182;
razn_w_mem[13359] = 182;
razn_w_mem[13360] = 182;
razn_w_mem[13361] = 182;
razn_w_mem[13362] = 182;
razn_w_mem[13363] = 182;
razn_w_mem[13364] = 182;
razn_w_mem[13365] = 182;
razn_w_mem[13366] = 182;
razn_w_mem[13367] = 182;
razn_w_mem[13368] = 182;
razn_w_mem[13369] = 182;
razn_w_mem[13370] = 182;
razn_w_mem[13371] = 182;
razn_w_mem[13372] = 182;
razn_w_mem[13373] = 182;
razn_w_mem[13374] = 182;
razn_w_mem[13375] = 182;
razn_w_mem[13376] = 182;
razn_w_mem[13377] = 182;
razn_w_mem[13378] = 182;
razn_w_mem[13379] = 182;
razn_w_mem[13380] = 182;
razn_w_mem[13381] = 182;
razn_w_mem[13382] = 182;
razn_w_mem[13383] = 182;
razn_w_mem[13384] = 182;
razn_w_mem[13385] = 182;
razn_w_mem[13386] = 182;
razn_w_mem[13387] = 182;
razn_w_mem[13388] = 182;
razn_w_mem[13389] = 182;
razn_w_mem[13390] = 182;
razn_w_mem[13391] = 182;
razn_w_mem[13392] = 182;
razn_w_mem[13393] = 182;
razn_w_mem[13394] = 182;
razn_w_mem[13395] = 182;
razn_w_mem[13396] = 182;
razn_w_mem[13397] = 182;
razn_w_mem[13398] = 182;
razn_w_mem[13399] = 182;
razn_w_mem[13400] = 182;
razn_w_mem[13401] = 182;
razn_w_mem[13402] = 182;
razn_w_mem[13403] = 182;
razn_w_mem[13404] = 182;
razn_w_mem[13405] = 182;
razn_w_mem[13406] = 182;
razn_w_mem[13407] = 182;
razn_w_mem[13408] = 182;
razn_w_mem[13409] = 182;
razn_w_mem[13410] = 182;
razn_w_mem[13411] = 182;
razn_w_mem[13412] = 182;
razn_w_mem[13413] = 182;
razn_w_mem[13414] = 182;
razn_w_mem[13415] = 182;
razn_w_mem[13416] = 182;
razn_w_mem[13417] = 182;
razn_w_mem[13418] = 182;
razn_w_mem[13419] = 182;
razn_w_mem[13420] = 182;
razn_w_mem[13421] = 182;
razn_w_mem[13422] = 182;
razn_w_mem[13423] = 182;
razn_w_mem[13424] = 182;
razn_w_mem[13425] = 182;
razn_w_mem[13426] = 182;
razn_w_mem[13427] = 182;
razn_w_mem[13428] = 182;
razn_w_mem[13429] = 182;
razn_w_mem[13430] = 182;
razn_w_mem[13431] = 182;
razn_w_mem[13432] = 182;
razn_w_mem[13433] = 182;
razn_w_mem[13434] = 182;
razn_w_mem[13435] = 182;
razn_w_mem[13436] = 182;
razn_w_mem[13437] = 182;
razn_w_mem[13438] = 182;
razn_w_mem[13439] = 182;
razn_w_mem[13440] = 152;
razn_w_mem[13441] = 152;
razn_w_mem[13442] = 152;
razn_w_mem[13443] = 152;
razn_w_mem[13444] = 152;
razn_w_mem[13445] = 152;
razn_w_mem[13446] = 152;
razn_w_mem[13447] = 152;
razn_w_mem[13448] = 152;
razn_w_mem[13449] = 152;
razn_w_mem[13450] = 152;
razn_w_mem[13451] = 152;
razn_w_mem[13452] = 152;
razn_w_mem[13453] = 152;
razn_w_mem[13454] = 152;
razn_w_mem[13455] = 152;
razn_w_mem[13456] = 152;
razn_w_mem[13457] = 152;
razn_w_mem[13458] = 152;
razn_w_mem[13459] = 152;
razn_w_mem[13460] = 152;
razn_w_mem[13461] = 152;
razn_w_mem[13462] = 152;
razn_w_mem[13463] = 152;
razn_w_mem[13464] = 152;
razn_w_mem[13465] = 152;
razn_w_mem[13466] = 152;
razn_w_mem[13467] = 152;
razn_w_mem[13468] = 152;
razn_w_mem[13469] = 152;
razn_w_mem[13470] = 152;
razn_w_mem[13471] = 152;
razn_w_mem[13472] = 152;
razn_w_mem[13473] = 152;
razn_w_mem[13474] = 152;
razn_w_mem[13475] = 152;
razn_w_mem[13476] = 152;
razn_w_mem[13477] = 152;
razn_w_mem[13478] = 152;
razn_w_mem[13479] = 152;
razn_w_mem[13480] = 152;
razn_w_mem[13481] = 152;
razn_w_mem[13482] = 152;
razn_w_mem[13483] = 152;
razn_w_mem[13484] = 152;
razn_w_mem[13485] = 152;
razn_w_mem[13486] = 152;
razn_w_mem[13487] = 152;
razn_w_mem[13488] = 152;
razn_w_mem[13489] = 152;
razn_w_mem[13490] = 152;
razn_w_mem[13491] = 152;
razn_w_mem[13492] = 152;
razn_w_mem[13493] = 152;
razn_w_mem[13494] = 152;
razn_w_mem[13495] = 152;
razn_w_mem[13496] = 152;
razn_w_mem[13497] = 152;
razn_w_mem[13498] = 152;
razn_w_mem[13499] = 152;
razn_w_mem[13500] = 152;
razn_w_mem[13501] = 152;
razn_w_mem[13502] = 152;
razn_w_mem[13503] = 152;
razn_w_mem[13504] = 152;
razn_w_mem[13505] = 152;
razn_w_mem[13506] = 152;
razn_w_mem[13507] = 152;
razn_w_mem[13508] = 152;
razn_w_mem[13509] = 152;
razn_w_mem[13510] = 152;
razn_w_mem[13511] = 152;
razn_w_mem[13512] = 152;
razn_w_mem[13513] = 152;
razn_w_mem[13514] = 152;
razn_w_mem[13515] = 152;
razn_w_mem[13516] = 152;
razn_w_mem[13517] = 152;
razn_w_mem[13518] = 152;
razn_w_mem[13519] = 152;
razn_w_mem[13520] = 152;
razn_w_mem[13521] = 152;
razn_w_mem[13522] = 152;
razn_w_mem[13523] = 152;
razn_w_mem[13524] = 152;
razn_w_mem[13525] = 152;
razn_w_mem[13526] = 152;
razn_w_mem[13527] = 152;
razn_w_mem[13528] = 152;
razn_w_mem[13529] = 152;
razn_w_mem[13530] = 152;
razn_w_mem[13531] = 152;
razn_w_mem[13532] = 152;
razn_w_mem[13533] = 152;
razn_w_mem[13534] = 152;
razn_w_mem[13535] = 152;
razn_w_mem[13536] = 152;
razn_w_mem[13537] = 152;
razn_w_mem[13538] = 152;
razn_w_mem[13539] = 152;
razn_w_mem[13540] = 152;
razn_w_mem[13541] = 152;
razn_w_mem[13542] = 152;
razn_w_mem[13543] = 152;
razn_w_mem[13544] = 152;
razn_w_mem[13545] = 152;
razn_w_mem[13546] = 152;
razn_w_mem[13547] = 152;
razn_w_mem[13548] = 152;
razn_w_mem[13549] = 152;
razn_w_mem[13550] = 152;
razn_w_mem[13551] = 152;
razn_w_mem[13552] = 152;
razn_w_mem[13553] = 152;
razn_w_mem[13554] = 152;
razn_w_mem[13555] = 152;
razn_w_mem[13556] = 152;
razn_w_mem[13557] = 152;
razn_w_mem[13558] = 152;
razn_w_mem[13559] = 152;
razn_w_mem[13560] = 152;
razn_w_mem[13561] = 152;
razn_w_mem[13562] = 152;
razn_w_mem[13563] = 152;
razn_w_mem[13564] = 152;
razn_w_mem[13565] = 152;
razn_w_mem[13566] = 152;
razn_w_mem[13567] = 152;
razn_w_mem[13568] = 122;
razn_w_mem[13569] = 122;
razn_w_mem[13570] = 122;
razn_w_mem[13571] = 122;
razn_w_mem[13572] = 122;
razn_w_mem[13573] = 122;
razn_w_mem[13574] = 122;
razn_w_mem[13575] = 122;
razn_w_mem[13576] = 122;
razn_w_mem[13577] = 122;
razn_w_mem[13578] = 122;
razn_w_mem[13579] = 122;
razn_w_mem[13580] = 122;
razn_w_mem[13581] = 122;
razn_w_mem[13582] = 122;
razn_w_mem[13583] = 122;
razn_w_mem[13584] = 122;
razn_w_mem[13585] = 122;
razn_w_mem[13586] = 122;
razn_w_mem[13587] = 122;
razn_w_mem[13588] = 122;
razn_w_mem[13589] = 122;
razn_w_mem[13590] = 122;
razn_w_mem[13591] = 122;
razn_w_mem[13592] = 122;
razn_w_mem[13593] = 122;
razn_w_mem[13594] = 122;
razn_w_mem[13595] = 122;
razn_w_mem[13596] = 122;
razn_w_mem[13597] = 122;
razn_w_mem[13598] = 122;
razn_w_mem[13599] = 122;
razn_w_mem[13600] = 122;
razn_w_mem[13601] = 122;
razn_w_mem[13602] = 122;
razn_w_mem[13603] = 122;
razn_w_mem[13604] = 122;
razn_w_mem[13605] = 122;
razn_w_mem[13606] = 122;
razn_w_mem[13607] = 122;
razn_w_mem[13608] = 122;
razn_w_mem[13609] = 122;
razn_w_mem[13610] = 122;
razn_w_mem[13611] = 122;
razn_w_mem[13612] = 122;
razn_w_mem[13613] = 122;
razn_w_mem[13614] = 122;
razn_w_mem[13615] = 122;
razn_w_mem[13616] = 122;
razn_w_mem[13617] = 122;
razn_w_mem[13618] = 122;
razn_w_mem[13619] = 122;
razn_w_mem[13620] = 122;
razn_w_mem[13621] = 122;
razn_w_mem[13622] = 122;
razn_w_mem[13623] = 122;
razn_w_mem[13624] = 122;
razn_w_mem[13625] = 122;
razn_w_mem[13626] = 122;
razn_w_mem[13627] = 122;
razn_w_mem[13628] = 122;
razn_w_mem[13629] = 122;
razn_w_mem[13630] = 122;
razn_w_mem[13631] = 122;
razn_w_mem[13632] = 122;
razn_w_mem[13633] = 122;
razn_w_mem[13634] = 122;
razn_w_mem[13635] = 122;
razn_w_mem[13636] = 122;
razn_w_mem[13637] = 122;
razn_w_mem[13638] = 122;
razn_w_mem[13639] = 122;
razn_w_mem[13640] = 122;
razn_w_mem[13641] = 122;
razn_w_mem[13642] = 122;
razn_w_mem[13643] = 122;
razn_w_mem[13644] = 122;
razn_w_mem[13645] = 122;
razn_w_mem[13646] = 122;
razn_w_mem[13647] = 122;
razn_w_mem[13648] = 122;
razn_w_mem[13649] = 122;
razn_w_mem[13650] = 122;
razn_w_mem[13651] = 122;
razn_w_mem[13652] = 122;
razn_w_mem[13653] = 122;
razn_w_mem[13654] = 122;
razn_w_mem[13655] = 122;
razn_w_mem[13656] = 122;
razn_w_mem[13657] = 122;
razn_w_mem[13658] = 122;
razn_w_mem[13659] = 122;
razn_w_mem[13660] = 122;
razn_w_mem[13661] = 122;
razn_w_mem[13662] = 122;
razn_w_mem[13663] = 122;
razn_w_mem[13664] = 122;
razn_w_mem[13665] = 122;
razn_w_mem[13666] = 122;
razn_w_mem[13667] = 122;
razn_w_mem[13668] = 122;
razn_w_mem[13669] = 122;
razn_w_mem[13670] = 122;
razn_w_mem[13671] = 122;
razn_w_mem[13672] = 122;
razn_w_mem[13673] = 122;
razn_w_mem[13674] = 122;
razn_w_mem[13675] = 122;
razn_w_mem[13676] = 122;
razn_w_mem[13677] = 122;
razn_w_mem[13678] = 122;
razn_w_mem[13679] = 122;
razn_w_mem[13680] = 122;
razn_w_mem[13681] = 122;
razn_w_mem[13682] = 122;
razn_w_mem[13683] = 122;
razn_w_mem[13684] = 122;
razn_w_mem[13685] = 122;
razn_w_mem[13686] = 122;
razn_w_mem[13687] = 122;
razn_w_mem[13688] = 122;
razn_w_mem[13689] = 122;
razn_w_mem[13690] = 122;
razn_w_mem[13691] = 122;
razn_w_mem[13692] = 122;
razn_w_mem[13693] = 122;
razn_w_mem[13694] = 122;
razn_w_mem[13695] = 122;
razn_w_mem[13696] = 92;
razn_w_mem[13697] = 92;
razn_w_mem[13698] = 92;
razn_w_mem[13699] = 92;
razn_w_mem[13700] = 92;
razn_w_mem[13701] = 92;
razn_w_mem[13702] = 92;
razn_w_mem[13703] = 92;
razn_w_mem[13704] = 92;
razn_w_mem[13705] = 92;
razn_w_mem[13706] = 92;
razn_w_mem[13707] = 92;
razn_w_mem[13708] = 92;
razn_w_mem[13709] = 92;
razn_w_mem[13710] = 92;
razn_w_mem[13711] = 92;
razn_w_mem[13712] = 92;
razn_w_mem[13713] = 92;
razn_w_mem[13714] = 92;
razn_w_mem[13715] = 92;
razn_w_mem[13716] = 92;
razn_w_mem[13717] = 92;
razn_w_mem[13718] = 92;
razn_w_mem[13719] = 92;
razn_w_mem[13720] = 92;
razn_w_mem[13721] = 92;
razn_w_mem[13722] = 92;
razn_w_mem[13723] = 92;
razn_w_mem[13724] = 92;
razn_w_mem[13725] = 92;
razn_w_mem[13726] = 92;
razn_w_mem[13727] = 92;
razn_w_mem[13728] = 92;
razn_w_mem[13729] = 92;
razn_w_mem[13730] = 92;
razn_w_mem[13731] = 92;
razn_w_mem[13732] = 92;
razn_w_mem[13733] = 92;
razn_w_mem[13734] = 92;
razn_w_mem[13735] = 92;
razn_w_mem[13736] = 92;
razn_w_mem[13737] = 92;
razn_w_mem[13738] = 92;
razn_w_mem[13739] = 92;
razn_w_mem[13740] = 92;
razn_w_mem[13741] = 92;
razn_w_mem[13742] = 92;
razn_w_mem[13743] = 92;
razn_w_mem[13744] = 92;
razn_w_mem[13745] = 92;
razn_w_mem[13746] = 92;
razn_w_mem[13747] = 92;
razn_w_mem[13748] = 92;
razn_w_mem[13749] = 92;
razn_w_mem[13750] = 92;
razn_w_mem[13751] = 92;
razn_w_mem[13752] = 92;
razn_w_mem[13753] = 92;
razn_w_mem[13754] = 92;
razn_w_mem[13755] = 92;
razn_w_mem[13756] = 92;
razn_w_mem[13757] = 92;
razn_w_mem[13758] = 92;
razn_w_mem[13759] = 92;
razn_w_mem[13760] = 92;
razn_w_mem[13761] = 92;
razn_w_mem[13762] = 92;
razn_w_mem[13763] = 92;
razn_w_mem[13764] = 92;
razn_w_mem[13765] = 92;
razn_w_mem[13766] = 92;
razn_w_mem[13767] = 92;
razn_w_mem[13768] = 92;
razn_w_mem[13769] = 92;
razn_w_mem[13770] = 92;
razn_w_mem[13771] = 92;
razn_w_mem[13772] = 92;
razn_w_mem[13773] = 92;
razn_w_mem[13774] = 92;
razn_w_mem[13775] = 92;
razn_w_mem[13776] = 92;
razn_w_mem[13777] = 92;
razn_w_mem[13778] = 92;
razn_w_mem[13779] = 92;
razn_w_mem[13780] = 92;
razn_w_mem[13781] = 92;
razn_w_mem[13782] = 92;
razn_w_mem[13783] = 92;
razn_w_mem[13784] = 92;
razn_w_mem[13785] = 92;
razn_w_mem[13786] = 92;
razn_w_mem[13787] = 92;
razn_w_mem[13788] = 92;
razn_w_mem[13789] = 92;
razn_w_mem[13790] = 92;
razn_w_mem[13791] = 92;
razn_w_mem[13792] = 92;
razn_w_mem[13793] = 92;
razn_w_mem[13794] = 92;
razn_w_mem[13795] = 92;
razn_w_mem[13796] = 92;
razn_w_mem[13797] = 92;
razn_w_mem[13798] = 92;
razn_w_mem[13799] = 92;
razn_w_mem[13800] = 92;
razn_w_mem[13801] = 92;
razn_w_mem[13802] = 92;
razn_w_mem[13803] = 92;
razn_w_mem[13804] = 92;
razn_w_mem[13805] = 92;
razn_w_mem[13806] = 92;
razn_w_mem[13807] = 92;
razn_w_mem[13808] = 92;
razn_w_mem[13809] = 92;
razn_w_mem[13810] = 92;
razn_w_mem[13811] = 92;
razn_w_mem[13812] = 92;
razn_w_mem[13813] = 92;
razn_w_mem[13814] = 92;
razn_w_mem[13815] = 92;
razn_w_mem[13816] = 92;
razn_w_mem[13817] = 92;
razn_w_mem[13818] = 92;
razn_w_mem[13819] = 92;
razn_w_mem[13820] = 92;
razn_w_mem[13821] = 92;
razn_w_mem[13822] = 92;
razn_w_mem[13823] = 92;
razn_w_mem[13824] = 62;
razn_w_mem[13825] = 62;
razn_w_mem[13826] = 62;
razn_w_mem[13827] = 62;
razn_w_mem[13828] = 62;
razn_w_mem[13829] = 62;
razn_w_mem[13830] = 62;
razn_w_mem[13831] = 62;
razn_w_mem[13832] = 62;
razn_w_mem[13833] = 62;
razn_w_mem[13834] = 62;
razn_w_mem[13835] = 62;
razn_w_mem[13836] = 62;
razn_w_mem[13837] = 62;
razn_w_mem[13838] = 62;
razn_w_mem[13839] = 62;
razn_w_mem[13840] = 62;
razn_w_mem[13841] = 62;
razn_w_mem[13842] = 62;
razn_w_mem[13843] = 62;
razn_w_mem[13844] = 62;
razn_w_mem[13845] = 62;
razn_w_mem[13846] = 62;
razn_w_mem[13847] = 62;
razn_w_mem[13848] = 62;
razn_w_mem[13849] = 62;
razn_w_mem[13850] = 62;
razn_w_mem[13851] = 62;
razn_w_mem[13852] = 62;
razn_w_mem[13853] = 62;
razn_w_mem[13854] = 62;
razn_w_mem[13855] = 62;
razn_w_mem[13856] = 62;
razn_w_mem[13857] = 62;
razn_w_mem[13858] = 62;
razn_w_mem[13859] = 62;
razn_w_mem[13860] = 62;
razn_w_mem[13861] = 62;
razn_w_mem[13862] = 62;
razn_w_mem[13863] = 62;
razn_w_mem[13864] = 62;
razn_w_mem[13865] = 62;
razn_w_mem[13866] = 62;
razn_w_mem[13867] = 62;
razn_w_mem[13868] = 62;
razn_w_mem[13869] = 62;
razn_w_mem[13870] = 62;
razn_w_mem[13871] = 62;
razn_w_mem[13872] = 62;
razn_w_mem[13873] = 62;
razn_w_mem[13874] = 62;
razn_w_mem[13875] = 62;
razn_w_mem[13876] = 62;
razn_w_mem[13877] = 62;
razn_w_mem[13878] = 62;
razn_w_mem[13879] = 62;
razn_w_mem[13880] = 62;
razn_w_mem[13881] = 62;
razn_w_mem[13882] = 62;
razn_w_mem[13883] = 62;
razn_w_mem[13884] = 62;
razn_w_mem[13885] = 62;
razn_w_mem[13886] = 62;
razn_w_mem[13887] = 62;
razn_w_mem[13888] = 62;
razn_w_mem[13889] = 62;
razn_w_mem[13890] = 62;
razn_w_mem[13891] = 62;
razn_w_mem[13892] = 62;
razn_w_mem[13893] = 62;
razn_w_mem[13894] = 62;
razn_w_mem[13895] = 62;
razn_w_mem[13896] = 62;
razn_w_mem[13897] = 62;
razn_w_mem[13898] = 62;
razn_w_mem[13899] = 62;
razn_w_mem[13900] = 62;
razn_w_mem[13901] = 62;
razn_w_mem[13902] = 62;
razn_w_mem[13903] = 62;
razn_w_mem[13904] = 62;
razn_w_mem[13905] = 62;
razn_w_mem[13906] = 62;
razn_w_mem[13907] = 62;
razn_w_mem[13908] = 62;
razn_w_mem[13909] = 62;
razn_w_mem[13910] = 62;
razn_w_mem[13911] = 62;
razn_w_mem[13912] = 62;
razn_w_mem[13913] = 62;
razn_w_mem[13914] = 62;
razn_w_mem[13915] = 62;
razn_w_mem[13916] = 62;
razn_w_mem[13917] = 62;
razn_w_mem[13918] = 62;
razn_w_mem[13919] = 62;
razn_w_mem[13920] = 62;
razn_w_mem[13921] = 62;
razn_w_mem[13922] = 62;
razn_w_mem[13923] = 62;
razn_w_mem[13924] = 62;
razn_w_mem[13925] = 62;
razn_w_mem[13926] = 62;
razn_w_mem[13927] = 62;
razn_w_mem[13928] = 62;
razn_w_mem[13929] = 62;
razn_w_mem[13930] = 62;
razn_w_mem[13931] = 62;
razn_w_mem[13932] = 62;
razn_w_mem[13933] = 62;
razn_w_mem[13934] = 62;
razn_w_mem[13935] = 62;
razn_w_mem[13936] = 62;
razn_w_mem[13937] = 62;
razn_w_mem[13938] = 62;
razn_w_mem[13939] = 62;
razn_w_mem[13940] = 62;
razn_w_mem[13941] = 62;
razn_w_mem[13942] = 62;
razn_w_mem[13943] = 62;
razn_w_mem[13944] = 62;
razn_w_mem[13945] = 62;
razn_w_mem[13946] = 62;
razn_w_mem[13947] = 62;
razn_w_mem[13948] = 62;
razn_w_mem[13949] = 62;
razn_w_mem[13950] = 62;
razn_w_mem[13951] = 62;
razn_w_mem[13952] = 32;
razn_w_mem[13953] = 32;
razn_w_mem[13954] = 32;
razn_w_mem[13955] = 32;
razn_w_mem[13956] = 32;
razn_w_mem[13957] = 32;
razn_w_mem[13958] = 32;
razn_w_mem[13959] = 32;
razn_w_mem[13960] = 32;
razn_w_mem[13961] = 32;
razn_w_mem[13962] = 32;
razn_w_mem[13963] = 32;
razn_w_mem[13964] = 32;
razn_w_mem[13965] = 32;
razn_w_mem[13966] = 32;
razn_w_mem[13967] = 32;
razn_w_mem[13968] = 32;
razn_w_mem[13969] = 32;
razn_w_mem[13970] = 32;
razn_w_mem[13971] = 32;
razn_w_mem[13972] = 32;
razn_w_mem[13973] = 32;
razn_w_mem[13974] = 32;
razn_w_mem[13975] = 32;
razn_w_mem[13976] = 32;
razn_w_mem[13977] = 32;
razn_w_mem[13978] = 32;
razn_w_mem[13979] = 32;
razn_w_mem[13980] = 32;
razn_w_mem[13981] = 32;
razn_w_mem[13982] = 32;
razn_w_mem[13983] = 32;
razn_w_mem[13984] = 32;
razn_w_mem[13985] = 32;
razn_w_mem[13986] = 32;
razn_w_mem[13987] = 32;
razn_w_mem[13988] = 32;
razn_w_mem[13989] = 32;
razn_w_mem[13990] = 32;
razn_w_mem[13991] = 32;
razn_w_mem[13992] = 32;
razn_w_mem[13993] = 32;
razn_w_mem[13994] = 32;
razn_w_mem[13995] = 32;
razn_w_mem[13996] = 32;
razn_w_mem[13997] = 32;
razn_w_mem[13998] = 32;
razn_w_mem[13999] = 32;
razn_w_mem[14000] = 32;
razn_w_mem[14001] = 32;
razn_w_mem[14002] = 32;
razn_w_mem[14003] = 32;
razn_w_mem[14004] = 32;
razn_w_mem[14005] = 32;
razn_w_mem[14006] = 32;
razn_w_mem[14007] = 32;
razn_w_mem[14008] = 32;
razn_w_mem[14009] = 32;
razn_w_mem[14010] = 32;
razn_w_mem[14011] = 32;
razn_w_mem[14012] = 32;
razn_w_mem[14013] = 32;
razn_w_mem[14014] = 32;
razn_w_mem[14015] = 32;
razn_w_mem[14016] = 32;
razn_w_mem[14017] = 32;
razn_w_mem[14018] = 32;
razn_w_mem[14019] = 32;
razn_w_mem[14020] = 32;
razn_w_mem[14021] = 32;
razn_w_mem[14022] = 32;
razn_w_mem[14023] = 32;
razn_w_mem[14024] = 32;
razn_w_mem[14025] = 32;
razn_w_mem[14026] = 32;
razn_w_mem[14027] = 32;
razn_w_mem[14028] = 32;
razn_w_mem[14029] = 32;
razn_w_mem[14030] = 32;
razn_w_mem[14031] = 32;
razn_w_mem[14032] = 32;
razn_w_mem[14033] = 32;
razn_w_mem[14034] = 32;
razn_w_mem[14035] = 32;
razn_w_mem[14036] = 32;
razn_w_mem[14037] = 32;
razn_w_mem[14038] = 32;
razn_w_mem[14039] = 32;
razn_w_mem[14040] = 32;
razn_w_mem[14041] = 32;
razn_w_mem[14042] = 32;
razn_w_mem[14043] = 32;
razn_w_mem[14044] = 32;
razn_w_mem[14045] = 32;
razn_w_mem[14046] = 32;
razn_w_mem[14047] = 32;
razn_w_mem[14048] = 32;
razn_w_mem[14049] = 32;
razn_w_mem[14050] = 32;
razn_w_mem[14051] = 32;
razn_w_mem[14052] = 32;
razn_w_mem[14053] = 32;
razn_w_mem[14054] = 32;
razn_w_mem[14055] = 32;
razn_w_mem[14056] = 32;
razn_w_mem[14057] = 32;
razn_w_mem[14058] = 32;
razn_w_mem[14059] = 32;
razn_w_mem[14060] = 32;
razn_w_mem[14061] = 32;
razn_w_mem[14062] = 32;
razn_w_mem[14063] = 32;
razn_w_mem[14064] = 32;
razn_w_mem[14065] = 32;
razn_w_mem[14066] = 32;
razn_w_mem[14067] = 32;
razn_w_mem[14068] = 32;
razn_w_mem[14069] = 32;
razn_w_mem[14070] = 32;
razn_w_mem[14071] = 32;
razn_w_mem[14072] = 32;
razn_w_mem[14073] = 32;
razn_w_mem[14074] = 32;
razn_w_mem[14075] = 32;
razn_w_mem[14076] = 32;
razn_w_mem[14077] = 32;
razn_w_mem[14078] = 32;
razn_w_mem[14079] = 32;
razn_w_mem[14080] = 2;
razn_w_mem[14081] = 2;
razn_w_mem[14082] = 2;
razn_w_mem[14083] = 2;
razn_w_mem[14084] = 2;
razn_w_mem[14085] = 2;
razn_w_mem[14086] = 2;
razn_w_mem[14087] = 2;
razn_w_mem[14088] = 2;
razn_w_mem[14089] = 2;
razn_w_mem[14090] = 2;
razn_w_mem[14091] = 2;
razn_w_mem[14092] = 2;
razn_w_mem[14093] = 2;
razn_w_mem[14094] = 2;
razn_w_mem[14095] = 2;
razn_w_mem[14096] = 2;
razn_w_mem[14097] = 2;
razn_w_mem[14098] = 2;
razn_w_mem[14099] = 2;
razn_w_mem[14100] = 2;
razn_w_mem[14101] = 2;
razn_w_mem[14102] = 2;
razn_w_mem[14103] = 2;
razn_w_mem[14104] = 2;
razn_w_mem[14105] = 2;
razn_w_mem[14106] = 2;
razn_w_mem[14107] = 2;
razn_w_mem[14108] = 2;
razn_w_mem[14109] = 2;
razn_w_mem[14110] = 2;
razn_w_mem[14111] = 2;
razn_w_mem[14112] = 2;
razn_w_mem[14113] = 2;
razn_w_mem[14114] = 2;
razn_w_mem[14115] = 2;
razn_w_mem[14116] = 2;
razn_w_mem[14117] = 2;
razn_w_mem[14118] = 2;
razn_w_mem[14119] = 2;
razn_w_mem[14120] = 2;
razn_w_mem[14121] = 2;
razn_w_mem[14122] = 2;
razn_w_mem[14123] = 2;
razn_w_mem[14124] = 2;
razn_w_mem[14125] = 2;
razn_w_mem[14126] = 2;
razn_w_mem[14127] = 2;
razn_w_mem[14128] = 2;
razn_w_mem[14129] = 2;
razn_w_mem[14130] = 2;
razn_w_mem[14131] = 2;
razn_w_mem[14132] = 2;
razn_w_mem[14133] = 2;
razn_w_mem[14134] = 2;
razn_w_mem[14135] = 2;
razn_w_mem[14136] = 2;
razn_w_mem[14137] = 2;
razn_w_mem[14138] = 2;
razn_w_mem[14139] = 2;
razn_w_mem[14140] = 2;
razn_w_mem[14141] = 2;
razn_w_mem[14142] = 2;
razn_w_mem[14143] = 2;
razn_w_mem[14144] = 2;
razn_w_mem[14145] = 2;
razn_w_mem[14146] = 2;
razn_w_mem[14147] = 2;
razn_w_mem[14148] = 2;
razn_w_mem[14149] = 2;
razn_w_mem[14150] = 2;
razn_w_mem[14151] = 2;
razn_w_mem[14152] = 2;
razn_w_mem[14153] = 2;
razn_w_mem[14154] = 2;
razn_w_mem[14155] = 2;
razn_w_mem[14156] = 2;
razn_w_mem[14157] = 2;
razn_w_mem[14158] = 2;
razn_w_mem[14159] = 2;
razn_w_mem[14160] = 2;
razn_w_mem[14161] = 2;
razn_w_mem[14162] = 2;
razn_w_mem[14163] = 2;
razn_w_mem[14164] = 2;
razn_w_mem[14165] = 2;
razn_w_mem[14166] = 2;
razn_w_mem[14167] = 2;
razn_w_mem[14168] = 2;
razn_w_mem[14169] = 2;
razn_w_mem[14170] = 2;
razn_w_mem[14171] = 2;
razn_w_mem[14172] = 2;
razn_w_mem[14173] = 2;
razn_w_mem[14174] = 2;
razn_w_mem[14175] = 2;
razn_w_mem[14176] = 2;
razn_w_mem[14177] = 2;
razn_w_mem[14178] = 2;
razn_w_mem[14179] = 2;
razn_w_mem[14180] = 2;
razn_w_mem[14181] = 2;
razn_w_mem[14182] = 2;
razn_w_mem[14183] = 2;
razn_w_mem[14184] = 2;
razn_w_mem[14185] = 2;
razn_w_mem[14186] = 2;
razn_w_mem[14187] = 2;
razn_w_mem[14188] = 2;
razn_w_mem[14189] = 2;
razn_w_mem[14190] = 2;
razn_w_mem[14191] = 2;
razn_w_mem[14192] = 2;
razn_w_mem[14193] = 2;
razn_w_mem[14194] = 2;
razn_w_mem[14195] = 2;
razn_w_mem[14196] = 2;
razn_w_mem[14197] = 2;
razn_w_mem[14198] = 2;
razn_w_mem[14199] = 2;
razn_w_mem[14200] = 2;
razn_w_mem[14201] = 2;
razn_w_mem[14202] = 2;
razn_w_mem[14203] = 2;
razn_w_mem[14204] = 2;
razn_w_mem[14205] = 2;
razn_w_mem[14206] = 2;
razn_w_mem[14207] = 2;
razn_w_mem[14208] = 226;
razn_w_mem[14209] = 226;
razn_w_mem[14210] = 226;
razn_w_mem[14211] = 226;
razn_w_mem[14212] = 226;
razn_w_mem[14213] = 226;
razn_w_mem[14214] = 226;
razn_w_mem[14215] = 226;
razn_w_mem[14216] = 226;
razn_w_mem[14217] = 226;
razn_w_mem[14218] = 226;
razn_w_mem[14219] = 226;
razn_w_mem[14220] = 226;
razn_w_mem[14221] = 226;
razn_w_mem[14222] = 226;
razn_w_mem[14223] = 226;
razn_w_mem[14224] = 226;
razn_w_mem[14225] = 226;
razn_w_mem[14226] = 226;
razn_w_mem[14227] = 226;
razn_w_mem[14228] = 226;
razn_w_mem[14229] = 226;
razn_w_mem[14230] = 226;
razn_w_mem[14231] = 226;
razn_w_mem[14232] = 226;
razn_w_mem[14233] = 226;
razn_w_mem[14234] = 226;
razn_w_mem[14235] = 226;
razn_w_mem[14236] = 226;
razn_w_mem[14237] = 226;
razn_w_mem[14238] = 226;
razn_w_mem[14239] = 226;
razn_w_mem[14240] = 226;
razn_w_mem[14241] = 226;
razn_w_mem[14242] = 226;
razn_w_mem[14243] = 226;
razn_w_mem[14244] = 226;
razn_w_mem[14245] = 226;
razn_w_mem[14246] = 226;
razn_w_mem[14247] = 226;
razn_w_mem[14248] = 226;
razn_w_mem[14249] = 226;
razn_w_mem[14250] = 226;
razn_w_mem[14251] = 226;
razn_w_mem[14252] = 226;
razn_w_mem[14253] = 226;
razn_w_mem[14254] = 226;
razn_w_mem[14255] = 226;
razn_w_mem[14256] = 226;
razn_w_mem[14257] = 226;
razn_w_mem[14258] = 226;
razn_w_mem[14259] = 226;
razn_w_mem[14260] = 226;
razn_w_mem[14261] = 226;
razn_w_mem[14262] = 226;
razn_w_mem[14263] = 226;
razn_w_mem[14264] = 226;
razn_w_mem[14265] = 226;
razn_w_mem[14266] = 226;
razn_w_mem[14267] = 226;
razn_w_mem[14268] = 226;
razn_w_mem[14269] = 226;
razn_w_mem[14270] = 226;
razn_w_mem[14271] = 226;
razn_w_mem[14272] = 226;
razn_w_mem[14273] = 226;
razn_w_mem[14274] = 226;
razn_w_mem[14275] = 226;
razn_w_mem[14276] = 226;
razn_w_mem[14277] = 226;
razn_w_mem[14278] = 226;
razn_w_mem[14279] = 226;
razn_w_mem[14280] = 226;
razn_w_mem[14281] = 226;
razn_w_mem[14282] = 226;
razn_w_mem[14283] = 226;
razn_w_mem[14284] = 226;
razn_w_mem[14285] = 226;
razn_w_mem[14286] = 226;
razn_w_mem[14287] = 226;
razn_w_mem[14288] = 226;
razn_w_mem[14289] = 226;
razn_w_mem[14290] = 226;
razn_w_mem[14291] = 226;
razn_w_mem[14292] = 226;
razn_w_mem[14293] = 226;
razn_w_mem[14294] = 226;
razn_w_mem[14295] = 226;
razn_w_mem[14296] = 226;
razn_w_mem[14297] = 226;
razn_w_mem[14298] = 226;
razn_w_mem[14299] = 226;
razn_w_mem[14300] = 226;
razn_w_mem[14301] = 226;
razn_w_mem[14302] = 226;
razn_w_mem[14303] = 226;
razn_w_mem[14304] = 226;
razn_w_mem[14305] = 226;
razn_w_mem[14306] = 226;
razn_w_mem[14307] = 226;
razn_w_mem[14308] = 226;
razn_w_mem[14309] = 226;
razn_w_mem[14310] = 226;
razn_w_mem[14311] = 226;
razn_w_mem[14312] = 226;
razn_w_mem[14313] = 226;
razn_w_mem[14314] = 226;
razn_w_mem[14315] = 226;
razn_w_mem[14316] = 226;
razn_w_mem[14317] = 226;
razn_w_mem[14318] = 226;
razn_w_mem[14319] = 226;
razn_w_mem[14320] = 226;
razn_w_mem[14321] = 226;
razn_w_mem[14322] = 226;
razn_w_mem[14323] = 226;
razn_w_mem[14324] = 226;
razn_w_mem[14325] = 226;
razn_w_mem[14326] = 226;
razn_w_mem[14327] = 226;
razn_w_mem[14328] = 226;
razn_w_mem[14329] = 226;
razn_w_mem[14330] = 226;
razn_w_mem[14331] = 226;
razn_w_mem[14332] = 226;
razn_w_mem[14333] = 226;
razn_w_mem[14334] = 226;
razn_w_mem[14335] = 226;
razn_w_mem[14336] = 196;
razn_w_mem[14337] = 196;
razn_w_mem[14338] = 196;
razn_w_mem[14339] = 196;
razn_w_mem[14340] = 196;
razn_w_mem[14341] = 196;
razn_w_mem[14342] = 196;
razn_w_mem[14343] = 196;
razn_w_mem[14344] = 196;
razn_w_mem[14345] = 196;
razn_w_mem[14346] = 196;
razn_w_mem[14347] = 196;
razn_w_mem[14348] = 196;
razn_w_mem[14349] = 196;
razn_w_mem[14350] = 196;
razn_w_mem[14351] = 196;
razn_w_mem[14352] = 196;
razn_w_mem[14353] = 196;
razn_w_mem[14354] = 196;
razn_w_mem[14355] = 196;
razn_w_mem[14356] = 196;
razn_w_mem[14357] = 196;
razn_w_mem[14358] = 196;
razn_w_mem[14359] = 196;
razn_w_mem[14360] = 196;
razn_w_mem[14361] = 196;
razn_w_mem[14362] = 196;
razn_w_mem[14363] = 196;
razn_w_mem[14364] = 196;
razn_w_mem[14365] = 196;
razn_w_mem[14366] = 196;
razn_w_mem[14367] = 196;
razn_w_mem[14368] = 196;
razn_w_mem[14369] = 196;
razn_w_mem[14370] = 196;
razn_w_mem[14371] = 196;
razn_w_mem[14372] = 196;
razn_w_mem[14373] = 196;
razn_w_mem[14374] = 196;
razn_w_mem[14375] = 196;
razn_w_mem[14376] = 196;
razn_w_mem[14377] = 196;
razn_w_mem[14378] = 196;
razn_w_mem[14379] = 196;
razn_w_mem[14380] = 196;
razn_w_mem[14381] = 196;
razn_w_mem[14382] = 196;
razn_w_mem[14383] = 196;
razn_w_mem[14384] = 196;
razn_w_mem[14385] = 196;
razn_w_mem[14386] = 196;
razn_w_mem[14387] = 196;
razn_w_mem[14388] = 196;
razn_w_mem[14389] = 196;
razn_w_mem[14390] = 196;
razn_w_mem[14391] = 196;
razn_w_mem[14392] = 196;
razn_w_mem[14393] = 196;
razn_w_mem[14394] = 196;
razn_w_mem[14395] = 196;
razn_w_mem[14396] = 196;
razn_w_mem[14397] = 196;
razn_w_mem[14398] = 196;
razn_w_mem[14399] = 196;
razn_w_mem[14400] = 196;
razn_w_mem[14401] = 196;
razn_w_mem[14402] = 196;
razn_w_mem[14403] = 196;
razn_w_mem[14404] = 196;
razn_w_mem[14405] = 196;
razn_w_mem[14406] = 196;
razn_w_mem[14407] = 196;
razn_w_mem[14408] = 196;
razn_w_mem[14409] = 196;
razn_w_mem[14410] = 196;
razn_w_mem[14411] = 196;
razn_w_mem[14412] = 196;
razn_w_mem[14413] = 196;
razn_w_mem[14414] = 196;
razn_w_mem[14415] = 196;
razn_w_mem[14416] = 196;
razn_w_mem[14417] = 196;
razn_w_mem[14418] = 196;
razn_w_mem[14419] = 196;
razn_w_mem[14420] = 196;
razn_w_mem[14421] = 196;
razn_w_mem[14422] = 196;
razn_w_mem[14423] = 196;
razn_w_mem[14424] = 196;
razn_w_mem[14425] = 196;
razn_w_mem[14426] = 196;
razn_w_mem[14427] = 196;
razn_w_mem[14428] = 196;
razn_w_mem[14429] = 196;
razn_w_mem[14430] = 196;
razn_w_mem[14431] = 196;
razn_w_mem[14432] = 196;
razn_w_mem[14433] = 196;
razn_w_mem[14434] = 196;
razn_w_mem[14435] = 196;
razn_w_mem[14436] = 196;
razn_w_mem[14437] = 196;
razn_w_mem[14438] = 196;
razn_w_mem[14439] = 196;
razn_w_mem[14440] = 196;
razn_w_mem[14441] = 196;
razn_w_mem[14442] = 196;
razn_w_mem[14443] = 196;
razn_w_mem[14444] = 196;
razn_w_mem[14445] = 196;
razn_w_mem[14446] = 196;
razn_w_mem[14447] = 196;
razn_w_mem[14448] = 196;
razn_w_mem[14449] = 196;
razn_w_mem[14450] = 196;
razn_w_mem[14451] = 196;
razn_w_mem[14452] = 196;
razn_w_mem[14453] = 196;
razn_w_mem[14454] = 196;
razn_w_mem[14455] = 196;
razn_w_mem[14456] = 196;
razn_w_mem[14457] = 196;
razn_w_mem[14458] = 196;
razn_w_mem[14459] = 196;
razn_w_mem[14460] = 196;
razn_w_mem[14461] = 196;
razn_w_mem[14462] = 196;
razn_w_mem[14463] = 196;
razn_w_mem[14464] = 166;
razn_w_mem[14465] = 166;
razn_w_mem[14466] = 166;
razn_w_mem[14467] = 166;
razn_w_mem[14468] = 166;
razn_w_mem[14469] = 166;
razn_w_mem[14470] = 166;
razn_w_mem[14471] = 166;
razn_w_mem[14472] = 166;
razn_w_mem[14473] = 166;
razn_w_mem[14474] = 166;
razn_w_mem[14475] = 166;
razn_w_mem[14476] = 166;
razn_w_mem[14477] = 166;
razn_w_mem[14478] = 166;
razn_w_mem[14479] = 166;
razn_w_mem[14480] = 166;
razn_w_mem[14481] = 166;
razn_w_mem[14482] = 166;
razn_w_mem[14483] = 166;
razn_w_mem[14484] = 166;
razn_w_mem[14485] = 166;
razn_w_mem[14486] = 166;
razn_w_mem[14487] = 166;
razn_w_mem[14488] = 166;
razn_w_mem[14489] = 166;
razn_w_mem[14490] = 166;
razn_w_mem[14491] = 166;
razn_w_mem[14492] = 166;
razn_w_mem[14493] = 166;
razn_w_mem[14494] = 166;
razn_w_mem[14495] = 166;
razn_w_mem[14496] = 166;
razn_w_mem[14497] = 166;
razn_w_mem[14498] = 166;
razn_w_mem[14499] = 166;
razn_w_mem[14500] = 166;
razn_w_mem[14501] = 166;
razn_w_mem[14502] = 166;
razn_w_mem[14503] = 166;
razn_w_mem[14504] = 166;
razn_w_mem[14505] = 166;
razn_w_mem[14506] = 166;
razn_w_mem[14507] = 166;
razn_w_mem[14508] = 166;
razn_w_mem[14509] = 166;
razn_w_mem[14510] = 166;
razn_w_mem[14511] = 166;
razn_w_mem[14512] = 166;
razn_w_mem[14513] = 166;
razn_w_mem[14514] = 166;
razn_w_mem[14515] = 166;
razn_w_mem[14516] = 166;
razn_w_mem[14517] = 166;
razn_w_mem[14518] = 166;
razn_w_mem[14519] = 166;
razn_w_mem[14520] = 166;
razn_w_mem[14521] = 166;
razn_w_mem[14522] = 166;
razn_w_mem[14523] = 166;
razn_w_mem[14524] = 166;
razn_w_mem[14525] = 166;
razn_w_mem[14526] = 166;
razn_w_mem[14527] = 166;
razn_w_mem[14528] = 166;
razn_w_mem[14529] = 166;
razn_w_mem[14530] = 166;
razn_w_mem[14531] = 166;
razn_w_mem[14532] = 166;
razn_w_mem[14533] = 166;
razn_w_mem[14534] = 166;
razn_w_mem[14535] = 166;
razn_w_mem[14536] = 166;
razn_w_mem[14537] = 166;
razn_w_mem[14538] = 166;
razn_w_mem[14539] = 166;
razn_w_mem[14540] = 166;
razn_w_mem[14541] = 166;
razn_w_mem[14542] = 166;
razn_w_mem[14543] = 166;
razn_w_mem[14544] = 166;
razn_w_mem[14545] = 166;
razn_w_mem[14546] = 166;
razn_w_mem[14547] = 166;
razn_w_mem[14548] = 166;
razn_w_mem[14549] = 166;
razn_w_mem[14550] = 166;
razn_w_mem[14551] = 166;
razn_w_mem[14552] = 166;
razn_w_mem[14553] = 166;
razn_w_mem[14554] = 166;
razn_w_mem[14555] = 166;
razn_w_mem[14556] = 166;
razn_w_mem[14557] = 166;
razn_w_mem[14558] = 166;
razn_w_mem[14559] = 166;
razn_w_mem[14560] = 166;
razn_w_mem[14561] = 166;
razn_w_mem[14562] = 166;
razn_w_mem[14563] = 166;
razn_w_mem[14564] = 166;
razn_w_mem[14565] = 166;
razn_w_mem[14566] = 166;
razn_w_mem[14567] = 166;
razn_w_mem[14568] = 166;
razn_w_mem[14569] = 166;
razn_w_mem[14570] = 166;
razn_w_mem[14571] = 166;
razn_w_mem[14572] = 166;
razn_w_mem[14573] = 166;
razn_w_mem[14574] = 166;
razn_w_mem[14575] = 166;
razn_w_mem[14576] = 166;
razn_w_mem[14577] = 166;
razn_w_mem[14578] = 166;
razn_w_mem[14579] = 166;
razn_w_mem[14580] = 166;
razn_w_mem[14581] = 166;
razn_w_mem[14582] = 166;
razn_w_mem[14583] = 166;
razn_w_mem[14584] = 166;
razn_w_mem[14585] = 166;
razn_w_mem[14586] = 166;
razn_w_mem[14587] = 166;
razn_w_mem[14588] = 166;
razn_w_mem[14589] = 166;
razn_w_mem[14590] = 166;
razn_w_mem[14591] = 166;
razn_w_mem[14592] = 136;
razn_w_mem[14593] = 136;
razn_w_mem[14594] = 136;
razn_w_mem[14595] = 136;
razn_w_mem[14596] = 136;
razn_w_mem[14597] = 136;
razn_w_mem[14598] = 136;
razn_w_mem[14599] = 136;
razn_w_mem[14600] = 136;
razn_w_mem[14601] = 136;
razn_w_mem[14602] = 136;
razn_w_mem[14603] = 136;
razn_w_mem[14604] = 136;
razn_w_mem[14605] = 136;
razn_w_mem[14606] = 136;
razn_w_mem[14607] = 136;
razn_w_mem[14608] = 136;
razn_w_mem[14609] = 136;
razn_w_mem[14610] = 136;
razn_w_mem[14611] = 136;
razn_w_mem[14612] = 136;
razn_w_mem[14613] = 136;
razn_w_mem[14614] = 136;
razn_w_mem[14615] = 136;
razn_w_mem[14616] = 136;
razn_w_mem[14617] = 136;
razn_w_mem[14618] = 136;
razn_w_mem[14619] = 136;
razn_w_mem[14620] = 136;
razn_w_mem[14621] = 136;
razn_w_mem[14622] = 136;
razn_w_mem[14623] = 136;
razn_w_mem[14624] = 136;
razn_w_mem[14625] = 136;
razn_w_mem[14626] = 136;
razn_w_mem[14627] = 136;
razn_w_mem[14628] = 136;
razn_w_mem[14629] = 136;
razn_w_mem[14630] = 136;
razn_w_mem[14631] = 136;
razn_w_mem[14632] = 136;
razn_w_mem[14633] = 136;
razn_w_mem[14634] = 136;
razn_w_mem[14635] = 136;
razn_w_mem[14636] = 136;
razn_w_mem[14637] = 136;
razn_w_mem[14638] = 136;
razn_w_mem[14639] = 136;
razn_w_mem[14640] = 136;
razn_w_mem[14641] = 136;
razn_w_mem[14642] = 136;
razn_w_mem[14643] = 136;
razn_w_mem[14644] = 136;
razn_w_mem[14645] = 136;
razn_w_mem[14646] = 136;
razn_w_mem[14647] = 136;
razn_w_mem[14648] = 136;
razn_w_mem[14649] = 136;
razn_w_mem[14650] = 136;
razn_w_mem[14651] = 136;
razn_w_mem[14652] = 136;
razn_w_mem[14653] = 136;
razn_w_mem[14654] = 136;
razn_w_mem[14655] = 136;
razn_w_mem[14656] = 136;
razn_w_mem[14657] = 136;
razn_w_mem[14658] = 136;
razn_w_mem[14659] = 136;
razn_w_mem[14660] = 136;
razn_w_mem[14661] = 136;
razn_w_mem[14662] = 136;
razn_w_mem[14663] = 136;
razn_w_mem[14664] = 136;
razn_w_mem[14665] = 136;
razn_w_mem[14666] = 136;
razn_w_mem[14667] = 136;
razn_w_mem[14668] = 136;
razn_w_mem[14669] = 136;
razn_w_mem[14670] = 136;
razn_w_mem[14671] = 136;
razn_w_mem[14672] = 136;
razn_w_mem[14673] = 136;
razn_w_mem[14674] = 136;
razn_w_mem[14675] = 136;
razn_w_mem[14676] = 136;
razn_w_mem[14677] = 136;
razn_w_mem[14678] = 136;
razn_w_mem[14679] = 136;
razn_w_mem[14680] = 136;
razn_w_mem[14681] = 136;
razn_w_mem[14682] = 136;
razn_w_mem[14683] = 136;
razn_w_mem[14684] = 136;
razn_w_mem[14685] = 136;
razn_w_mem[14686] = 136;
razn_w_mem[14687] = 136;
razn_w_mem[14688] = 136;
razn_w_mem[14689] = 136;
razn_w_mem[14690] = 136;
razn_w_mem[14691] = 136;
razn_w_mem[14692] = 136;
razn_w_mem[14693] = 136;
razn_w_mem[14694] = 136;
razn_w_mem[14695] = 136;
razn_w_mem[14696] = 136;
razn_w_mem[14697] = 136;
razn_w_mem[14698] = 136;
razn_w_mem[14699] = 136;
razn_w_mem[14700] = 136;
razn_w_mem[14701] = 136;
razn_w_mem[14702] = 136;
razn_w_mem[14703] = 136;
razn_w_mem[14704] = 136;
razn_w_mem[14705] = 136;
razn_w_mem[14706] = 136;
razn_w_mem[14707] = 136;
razn_w_mem[14708] = 136;
razn_w_mem[14709] = 136;
razn_w_mem[14710] = 136;
razn_w_mem[14711] = 136;
razn_w_mem[14712] = 136;
razn_w_mem[14713] = 136;
razn_w_mem[14714] = 136;
razn_w_mem[14715] = 136;
razn_w_mem[14716] = 136;
razn_w_mem[14717] = 136;
razn_w_mem[14718] = 136;
razn_w_mem[14719] = 136;
razn_w_mem[14720] = 106;
razn_w_mem[14721] = 106;
razn_w_mem[14722] = 106;
razn_w_mem[14723] = 106;
razn_w_mem[14724] = 106;
razn_w_mem[14725] = 106;
razn_w_mem[14726] = 106;
razn_w_mem[14727] = 106;
razn_w_mem[14728] = 106;
razn_w_mem[14729] = 106;
razn_w_mem[14730] = 106;
razn_w_mem[14731] = 106;
razn_w_mem[14732] = 106;
razn_w_mem[14733] = 106;
razn_w_mem[14734] = 106;
razn_w_mem[14735] = 106;
razn_w_mem[14736] = 106;
razn_w_mem[14737] = 106;
razn_w_mem[14738] = 106;
razn_w_mem[14739] = 106;
razn_w_mem[14740] = 106;
razn_w_mem[14741] = 106;
razn_w_mem[14742] = 106;
razn_w_mem[14743] = 106;
razn_w_mem[14744] = 106;
razn_w_mem[14745] = 106;
razn_w_mem[14746] = 106;
razn_w_mem[14747] = 106;
razn_w_mem[14748] = 106;
razn_w_mem[14749] = 106;
razn_w_mem[14750] = 106;
razn_w_mem[14751] = 106;
razn_w_mem[14752] = 106;
razn_w_mem[14753] = 106;
razn_w_mem[14754] = 106;
razn_w_mem[14755] = 106;
razn_w_mem[14756] = 106;
razn_w_mem[14757] = 106;
razn_w_mem[14758] = 106;
razn_w_mem[14759] = 106;
razn_w_mem[14760] = 106;
razn_w_mem[14761] = 106;
razn_w_mem[14762] = 106;
razn_w_mem[14763] = 106;
razn_w_mem[14764] = 106;
razn_w_mem[14765] = 106;
razn_w_mem[14766] = 106;
razn_w_mem[14767] = 106;
razn_w_mem[14768] = 106;
razn_w_mem[14769] = 106;
razn_w_mem[14770] = 106;
razn_w_mem[14771] = 106;
razn_w_mem[14772] = 106;
razn_w_mem[14773] = 106;
razn_w_mem[14774] = 106;
razn_w_mem[14775] = 106;
razn_w_mem[14776] = 106;
razn_w_mem[14777] = 106;
razn_w_mem[14778] = 106;
razn_w_mem[14779] = 106;
razn_w_mem[14780] = 106;
razn_w_mem[14781] = 106;
razn_w_mem[14782] = 106;
razn_w_mem[14783] = 106;
razn_w_mem[14784] = 106;
razn_w_mem[14785] = 106;
razn_w_mem[14786] = 106;
razn_w_mem[14787] = 106;
razn_w_mem[14788] = 106;
razn_w_mem[14789] = 106;
razn_w_mem[14790] = 106;
razn_w_mem[14791] = 106;
razn_w_mem[14792] = 106;
razn_w_mem[14793] = 106;
razn_w_mem[14794] = 106;
razn_w_mem[14795] = 106;
razn_w_mem[14796] = 106;
razn_w_mem[14797] = 106;
razn_w_mem[14798] = 106;
razn_w_mem[14799] = 106;
razn_w_mem[14800] = 106;
razn_w_mem[14801] = 106;
razn_w_mem[14802] = 106;
razn_w_mem[14803] = 106;
razn_w_mem[14804] = 106;
razn_w_mem[14805] = 106;
razn_w_mem[14806] = 106;
razn_w_mem[14807] = 106;
razn_w_mem[14808] = 106;
razn_w_mem[14809] = 106;
razn_w_mem[14810] = 106;
razn_w_mem[14811] = 106;
razn_w_mem[14812] = 106;
razn_w_mem[14813] = 106;
razn_w_mem[14814] = 106;
razn_w_mem[14815] = 106;
razn_w_mem[14816] = 106;
razn_w_mem[14817] = 106;
razn_w_mem[14818] = 106;
razn_w_mem[14819] = 106;
razn_w_mem[14820] = 106;
razn_w_mem[14821] = 106;
razn_w_mem[14822] = 106;
razn_w_mem[14823] = 106;
razn_w_mem[14824] = 106;
razn_w_mem[14825] = 106;
razn_w_mem[14826] = 106;
razn_w_mem[14827] = 106;
razn_w_mem[14828] = 106;
razn_w_mem[14829] = 106;
razn_w_mem[14830] = 106;
razn_w_mem[14831] = 106;
razn_w_mem[14832] = 106;
razn_w_mem[14833] = 106;
razn_w_mem[14834] = 106;
razn_w_mem[14835] = 106;
razn_w_mem[14836] = 106;
razn_w_mem[14837] = 106;
razn_w_mem[14838] = 106;
razn_w_mem[14839] = 106;
razn_w_mem[14840] = 106;
razn_w_mem[14841] = 106;
razn_w_mem[14842] = 106;
razn_w_mem[14843] = 106;
razn_w_mem[14844] = 106;
razn_w_mem[14845] = 106;
razn_w_mem[14846] = 106;
razn_w_mem[14847] = 106;
razn_w_mem[14848] = 76;
razn_w_mem[14849] = 76;
razn_w_mem[14850] = 76;
razn_w_mem[14851] = 76;
razn_w_mem[14852] = 76;
razn_w_mem[14853] = 76;
razn_w_mem[14854] = 76;
razn_w_mem[14855] = 76;
razn_w_mem[14856] = 76;
razn_w_mem[14857] = 76;
razn_w_mem[14858] = 76;
razn_w_mem[14859] = 76;
razn_w_mem[14860] = 76;
razn_w_mem[14861] = 76;
razn_w_mem[14862] = 76;
razn_w_mem[14863] = 76;
razn_w_mem[14864] = 76;
razn_w_mem[14865] = 76;
razn_w_mem[14866] = 76;
razn_w_mem[14867] = 76;
razn_w_mem[14868] = 76;
razn_w_mem[14869] = 76;
razn_w_mem[14870] = 76;
razn_w_mem[14871] = 76;
razn_w_mem[14872] = 76;
razn_w_mem[14873] = 76;
razn_w_mem[14874] = 76;
razn_w_mem[14875] = 76;
razn_w_mem[14876] = 76;
razn_w_mem[14877] = 76;
razn_w_mem[14878] = 76;
razn_w_mem[14879] = 76;
razn_w_mem[14880] = 76;
razn_w_mem[14881] = 76;
razn_w_mem[14882] = 76;
razn_w_mem[14883] = 76;
razn_w_mem[14884] = 76;
razn_w_mem[14885] = 76;
razn_w_mem[14886] = 76;
razn_w_mem[14887] = 76;
razn_w_mem[14888] = 76;
razn_w_mem[14889] = 76;
razn_w_mem[14890] = 76;
razn_w_mem[14891] = 76;
razn_w_mem[14892] = 76;
razn_w_mem[14893] = 76;
razn_w_mem[14894] = 76;
razn_w_mem[14895] = 76;
razn_w_mem[14896] = 76;
razn_w_mem[14897] = 76;
razn_w_mem[14898] = 76;
razn_w_mem[14899] = 76;
razn_w_mem[14900] = 76;
razn_w_mem[14901] = 76;
razn_w_mem[14902] = 76;
razn_w_mem[14903] = 76;
razn_w_mem[14904] = 76;
razn_w_mem[14905] = 76;
razn_w_mem[14906] = 76;
razn_w_mem[14907] = 76;
razn_w_mem[14908] = 76;
razn_w_mem[14909] = 76;
razn_w_mem[14910] = 76;
razn_w_mem[14911] = 76;
razn_w_mem[14912] = 76;
razn_w_mem[14913] = 76;
razn_w_mem[14914] = 76;
razn_w_mem[14915] = 76;
razn_w_mem[14916] = 76;
razn_w_mem[14917] = 76;
razn_w_mem[14918] = 76;
razn_w_mem[14919] = 76;
razn_w_mem[14920] = 76;
razn_w_mem[14921] = 76;
razn_w_mem[14922] = 76;
razn_w_mem[14923] = 76;
razn_w_mem[14924] = 76;
razn_w_mem[14925] = 76;
razn_w_mem[14926] = 76;
razn_w_mem[14927] = 76;
razn_w_mem[14928] = 76;
razn_w_mem[14929] = 76;
razn_w_mem[14930] = 76;
razn_w_mem[14931] = 76;
razn_w_mem[14932] = 76;
razn_w_mem[14933] = 76;
razn_w_mem[14934] = 76;
razn_w_mem[14935] = 76;
razn_w_mem[14936] = 76;
razn_w_mem[14937] = 76;
razn_w_mem[14938] = 76;
razn_w_mem[14939] = 76;
razn_w_mem[14940] = 76;
razn_w_mem[14941] = 76;
razn_w_mem[14942] = 76;
razn_w_mem[14943] = 76;
razn_w_mem[14944] = 76;
razn_w_mem[14945] = 76;
razn_w_mem[14946] = 76;
razn_w_mem[14947] = 76;
razn_w_mem[14948] = 76;
razn_w_mem[14949] = 76;
razn_w_mem[14950] = 76;
razn_w_mem[14951] = 76;
razn_w_mem[14952] = 76;
razn_w_mem[14953] = 76;
razn_w_mem[14954] = 76;
razn_w_mem[14955] = 76;
razn_w_mem[14956] = 76;
razn_w_mem[14957] = 76;
razn_w_mem[14958] = 76;
razn_w_mem[14959] = 76;
razn_w_mem[14960] = 76;
razn_w_mem[14961] = 76;
razn_w_mem[14962] = 76;
razn_w_mem[14963] = 76;
razn_w_mem[14964] = 76;
razn_w_mem[14965] = 76;
razn_w_mem[14966] = 76;
razn_w_mem[14967] = 76;
razn_w_mem[14968] = 76;
razn_w_mem[14969] = 76;
razn_w_mem[14970] = 76;
razn_w_mem[14971] = 76;
razn_w_mem[14972] = 76;
razn_w_mem[14973] = 76;
razn_w_mem[14974] = 76;
razn_w_mem[14975] = 76;
razn_w_mem[14976] = 46;
razn_w_mem[14977] = 46;
razn_w_mem[14978] = 46;
razn_w_mem[14979] = 46;
razn_w_mem[14980] = 46;
razn_w_mem[14981] = 46;
razn_w_mem[14982] = 46;
razn_w_mem[14983] = 46;
razn_w_mem[14984] = 46;
razn_w_mem[14985] = 46;
razn_w_mem[14986] = 46;
razn_w_mem[14987] = 46;
razn_w_mem[14988] = 46;
razn_w_mem[14989] = 46;
razn_w_mem[14990] = 46;
razn_w_mem[14991] = 46;
razn_w_mem[14992] = 46;
razn_w_mem[14993] = 46;
razn_w_mem[14994] = 46;
razn_w_mem[14995] = 46;
razn_w_mem[14996] = 46;
razn_w_mem[14997] = 46;
razn_w_mem[14998] = 46;
razn_w_mem[14999] = 46;
razn_w_mem[15000] = 46;
razn_w_mem[15001] = 46;
razn_w_mem[15002] = 46;
razn_w_mem[15003] = 46;
razn_w_mem[15004] = 46;
razn_w_mem[15005] = 46;
razn_w_mem[15006] = 46;
razn_w_mem[15007] = 46;
razn_w_mem[15008] = 46;
razn_w_mem[15009] = 46;
razn_w_mem[15010] = 46;
razn_w_mem[15011] = 46;
razn_w_mem[15012] = 46;
razn_w_mem[15013] = 46;
razn_w_mem[15014] = 46;
razn_w_mem[15015] = 46;
razn_w_mem[15016] = 46;
razn_w_mem[15017] = 46;
razn_w_mem[15018] = 46;
razn_w_mem[15019] = 46;
razn_w_mem[15020] = 46;
razn_w_mem[15021] = 46;
razn_w_mem[15022] = 46;
razn_w_mem[15023] = 46;
razn_w_mem[15024] = 46;
razn_w_mem[15025] = 46;
razn_w_mem[15026] = 46;
razn_w_mem[15027] = 46;
razn_w_mem[15028] = 46;
razn_w_mem[15029] = 46;
razn_w_mem[15030] = 46;
razn_w_mem[15031] = 46;
razn_w_mem[15032] = 46;
razn_w_mem[15033] = 46;
razn_w_mem[15034] = 46;
razn_w_mem[15035] = 46;
razn_w_mem[15036] = 46;
razn_w_mem[15037] = 46;
razn_w_mem[15038] = 46;
razn_w_mem[15039] = 46;
razn_w_mem[15040] = 46;
razn_w_mem[15041] = 46;
razn_w_mem[15042] = 46;
razn_w_mem[15043] = 46;
razn_w_mem[15044] = 46;
razn_w_mem[15045] = 46;
razn_w_mem[15046] = 46;
razn_w_mem[15047] = 46;
razn_w_mem[15048] = 46;
razn_w_mem[15049] = 46;
razn_w_mem[15050] = 46;
razn_w_mem[15051] = 46;
razn_w_mem[15052] = 46;
razn_w_mem[15053] = 46;
razn_w_mem[15054] = 46;
razn_w_mem[15055] = 46;
razn_w_mem[15056] = 46;
razn_w_mem[15057] = 46;
razn_w_mem[15058] = 46;
razn_w_mem[15059] = 46;
razn_w_mem[15060] = 46;
razn_w_mem[15061] = 46;
razn_w_mem[15062] = 46;
razn_w_mem[15063] = 46;
razn_w_mem[15064] = 46;
razn_w_mem[15065] = 46;
razn_w_mem[15066] = 46;
razn_w_mem[15067] = 46;
razn_w_mem[15068] = 46;
razn_w_mem[15069] = 46;
razn_w_mem[15070] = 46;
razn_w_mem[15071] = 46;
razn_w_mem[15072] = 46;
razn_w_mem[15073] = 46;
razn_w_mem[15074] = 46;
razn_w_mem[15075] = 46;
razn_w_mem[15076] = 46;
razn_w_mem[15077] = 46;
razn_w_mem[15078] = 46;
razn_w_mem[15079] = 46;
razn_w_mem[15080] = 46;
razn_w_mem[15081] = 46;
razn_w_mem[15082] = 46;
razn_w_mem[15083] = 46;
razn_w_mem[15084] = 46;
razn_w_mem[15085] = 46;
razn_w_mem[15086] = 46;
razn_w_mem[15087] = 46;
razn_w_mem[15088] = 46;
razn_w_mem[15089] = 46;
razn_w_mem[15090] = 46;
razn_w_mem[15091] = 46;
razn_w_mem[15092] = 46;
razn_w_mem[15093] = 46;
razn_w_mem[15094] = 46;
razn_w_mem[15095] = 46;
razn_w_mem[15096] = 46;
razn_w_mem[15097] = 46;
razn_w_mem[15098] = 46;
razn_w_mem[15099] = 46;
razn_w_mem[15100] = 46;
razn_w_mem[15101] = 46;
razn_w_mem[15102] = 46;
razn_w_mem[15103] = 46;
razn_w_mem[15104] = 16;
razn_w_mem[15105] = 16;
razn_w_mem[15106] = 16;
razn_w_mem[15107] = 16;
razn_w_mem[15108] = 16;
razn_w_mem[15109] = 16;
razn_w_mem[15110] = 16;
razn_w_mem[15111] = 16;
razn_w_mem[15112] = 16;
razn_w_mem[15113] = 16;
razn_w_mem[15114] = 16;
razn_w_mem[15115] = 16;
razn_w_mem[15116] = 16;
razn_w_mem[15117] = 16;
razn_w_mem[15118] = 16;
razn_w_mem[15119] = 16;
razn_w_mem[15120] = 16;
razn_w_mem[15121] = 16;
razn_w_mem[15122] = 16;
razn_w_mem[15123] = 16;
razn_w_mem[15124] = 16;
razn_w_mem[15125] = 16;
razn_w_mem[15126] = 16;
razn_w_mem[15127] = 16;
razn_w_mem[15128] = 16;
razn_w_mem[15129] = 16;
razn_w_mem[15130] = 16;
razn_w_mem[15131] = 16;
razn_w_mem[15132] = 16;
razn_w_mem[15133] = 16;
razn_w_mem[15134] = 16;
razn_w_mem[15135] = 16;
razn_w_mem[15136] = 16;
razn_w_mem[15137] = 16;
razn_w_mem[15138] = 16;
razn_w_mem[15139] = 16;
razn_w_mem[15140] = 16;
razn_w_mem[15141] = 16;
razn_w_mem[15142] = 16;
razn_w_mem[15143] = 16;
razn_w_mem[15144] = 16;
razn_w_mem[15145] = 16;
razn_w_mem[15146] = 16;
razn_w_mem[15147] = 16;
razn_w_mem[15148] = 16;
razn_w_mem[15149] = 16;
razn_w_mem[15150] = 16;
razn_w_mem[15151] = 16;
razn_w_mem[15152] = 16;
razn_w_mem[15153] = 16;
razn_w_mem[15154] = 16;
razn_w_mem[15155] = 16;
razn_w_mem[15156] = 16;
razn_w_mem[15157] = 16;
razn_w_mem[15158] = 16;
razn_w_mem[15159] = 16;
razn_w_mem[15160] = 16;
razn_w_mem[15161] = 16;
razn_w_mem[15162] = 16;
razn_w_mem[15163] = 16;
razn_w_mem[15164] = 16;
razn_w_mem[15165] = 16;
razn_w_mem[15166] = 16;
razn_w_mem[15167] = 16;
razn_w_mem[15168] = 16;
razn_w_mem[15169] = 16;
razn_w_mem[15170] = 16;
razn_w_mem[15171] = 16;
razn_w_mem[15172] = 16;
razn_w_mem[15173] = 16;
razn_w_mem[15174] = 16;
razn_w_mem[15175] = 16;
razn_w_mem[15176] = 16;
razn_w_mem[15177] = 16;
razn_w_mem[15178] = 16;
razn_w_mem[15179] = 16;
razn_w_mem[15180] = 16;
razn_w_mem[15181] = 16;
razn_w_mem[15182] = 16;
razn_w_mem[15183] = 16;
razn_w_mem[15184] = 16;
razn_w_mem[15185] = 16;
razn_w_mem[15186] = 16;
razn_w_mem[15187] = 16;
razn_w_mem[15188] = 16;
razn_w_mem[15189] = 16;
razn_w_mem[15190] = 16;
razn_w_mem[15191] = 16;
razn_w_mem[15192] = 16;
razn_w_mem[15193] = 16;
razn_w_mem[15194] = 16;
razn_w_mem[15195] = 16;
razn_w_mem[15196] = 16;
razn_w_mem[15197] = 16;
razn_w_mem[15198] = 16;
razn_w_mem[15199] = 16;
razn_w_mem[15200] = 16;
razn_w_mem[15201] = 16;
razn_w_mem[15202] = 16;
razn_w_mem[15203] = 16;
razn_w_mem[15204] = 16;
razn_w_mem[15205] = 16;
razn_w_mem[15206] = 16;
razn_w_mem[15207] = 16;
razn_w_mem[15208] = 16;
razn_w_mem[15209] = 16;
razn_w_mem[15210] = 16;
razn_w_mem[15211] = 16;
razn_w_mem[15212] = 16;
razn_w_mem[15213] = 16;
razn_w_mem[15214] = 16;
razn_w_mem[15215] = 16;
razn_w_mem[15216] = 16;
razn_w_mem[15217] = 16;
razn_w_mem[15218] = 16;
razn_w_mem[15219] = 16;
razn_w_mem[15220] = 16;
razn_w_mem[15221] = 16;
razn_w_mem[15222] = 16;
razn_w_mem[15223] = 16;
razn_w_mem[15224] = 16;
razn_w_mem[15225] = 16;
razn_w_mem[15226] = 16;
razn_w_mem[15227] = 16;
razn_w_mem[15228] = 16;
razn_w_mem[15229] = 16;
razn_w_mem[15230] = 16;
razn_w_mem[15231] = 16;
razn_w_mem[15232] = 240;
razn_w_mem[15233] = 240;
razn_w_mem[15234] = 240;
razn_w_mem[15235] = 240;
razn_w_mem[15236] = 240;
razn_w_mem[15237] = 240;
razn_w_mem[15238] = 240;
razn_w_mem[15239] = 240;
razn_w_mem[15240] = 240;
razn_w_mem[15241] = 240;
razn_w_mem[15242] = 240;
razn_w_mem[15243] = 240;
razn_w_mem[15244] = 240;
razn_w_mem[15245] = 240;
razn_w_mem[15246] = 240;
razn_w_mem[15247] = 240;
razn_w_mem[15248] = 240;
razn_w_mem[15249] = 240;
razn_w_mem[15250] = 240;
razn_w_mem[15251] = 240;
razn_w_mem[15252] = 240;
razn_w_mem[15253] = 240;
razn_w_mem[15254] = 240;
razn_w_mem[15255] = 240;
razn_w_mem[15256] = 240;
razn_w_mem[15257] = 240;
razn_w_mem[15258] = 240;
razn_w_mem[15259] = 240;
razn_w_mem[15260] = 240;
razn_w_mem[15261] = 240;
razn_w_mem[15262] = 240;
razn_w_mem[15263] = 240;
razn_w_mem[15264] = 240;
razn_w_mem[15265] = 240;
razn_w_mem[15266] = 240;
razn_w_mem[15267] = 240;
razn_w_mem[15268] = 240;
razn_w_mem[15269] = 240;
razn_w_mem[15270] = 240;
razn_w_mem[15271] = 240;
razn_w_mem[15272] = 240;
razn_w_mem[15273] = 240;
razn_w_mem[15274] = 240;
razn_w_mem[15275] = 240;
razn_w_mem[15276] = 240;
razn_w_mem[15277] = 240;
razn_w_mem[15278] = 240;
razn_w_mem[15279] = 240;
razn_w_mem[15280] = 240;
razn_w_mem[15281] = 240;
razn_w_mem[15282] = 240;
razn_w_mem[15283] = 240;
razn_w_mem[15284] = 240;
razn_w_mem[15285] = 240;
razn_w_mem[15286] = 240;
razn_w_mem[15287] = 240;
razn_w_mem[15288] = 240;
razn_w_mem[15289] = 240;
razn_w_mem[15290] = 240;
razn_w_mem[15291] = 240;
razn_w_mem[15292] = 240;
razn_w_mem[15293] = 240;
razn_w_mem[15294] = 240;
razn_w_mem[15295] = 240;
razn_w_mem[15296] = 240;
razn_w_mem[15297] = 240;
razn_w_mem[15298] = 240;
razn_w_mem[15299] = 240;
razn_w_mem[15300] = 240;
razn_w_mem[15301] = 240;
razn_w_mem[15302] = 240;
razn_w_mem[15303] = 240;
razn_w_mem[15304] = 240;
razn_w_mem[15305] = 240;
razn_w_mem[15306] = 240;
razn_w_mem[15307] = 240;
razn_w_mem[15308] = 240;
razn_w_mem[15309] = 240;
razn_w_mem[15310] = 240;
razn_w_mem[15311] = 240;
razn_w_mem[15312] = 240;
razn_w_mem[15313] = 240;
razn_w_mem[15314] = 240;
razn_w_mem[15315] = 240;
razn_w_mem[15316] = 240;
razn_w_mem[15317] = 240;
razn_w_mem[15318] = 240;
razn_w_mem[15319] = 240;
razn_w_mem[15320] = 240;
razn_w_mem[15321] = 240;
razn_w_mem[15322] = 240;
razn_w_mem[15323] = 240;
razn_w_mem[15324] = 240;
razn_w_mem[15325] = 240;
razn_w_mem[15326] = 240;
razn_w_mem[15327] = 240;
razn_w_mem[15328] = 240;
razn_w_mem[15329] = 240;
razn_w_mem[15330] = 240;
razn_w_mem[15331] = 240;
razn_w_mem[15332] = 240;
razn_w_mem[15333] = 240;
razn_w_mem[15334] = 240;
razn_w_mem[15335] = 240;
razn_w_mem[15336] = 240;
razn_w_mem[15337] = 240;
razn_w_mem[15338] = 240;
razn_w_mem[15339] = 240;
razn_w_mem[15340] = 240;
razn_w_mem[15341] = 240;
razn_w_mem[15342] = 240;
razn_w_mem[15343] = 240;
razn_w_mem[15344] = 240;
razn_w_mem[15345] = 240;
razn_w_mem[15346] = 240;
razn_w_mem[15347] = 240;
razn_w_mem[15348] = 240;
razn_w_mem[15349] = 240;
razn_w_mem[15350] = 240;
razn_w_mem[15351] = 240;
razn_w_mem[15352] = 240;
razn_w_mem[15353] = 240;
razn_w_mem[15354] = 240;
razn_w_mem[15355] = 240;
razn_w_mem[15356] = 240;
razn_w_mem[15357] = 240;
razn_w_mem[15358] = 240;
razn_w_mem[15359] = 240;
razn_w_mem[15360] = 210;
razn_w_mem[15361] = 210;
razn_w_mem[15362] = 210;
razn_w_mem[15363] = 210;
razn_w_mem[15364] = 210;
razn_w_mem[15365] = 210;
razn_w_mem[15366] = 210;
razn_w_mem[15367] = 210;
razn_w_mem[15368] = 210;
razn_w_mem[15369] = 210;
razn_w_mem[15370] = 210;
razn_w_mem[15371] = 210;
razn_w_mem[15372] = 210;
razn_w_mem[15373] = 210;
razn_w_mem[15374] = 210;
razn_w_mem[15375] = 210;
razn_w_mem[15376] = 210;
razn_w_mem[15377] = 210;
razn_w_mem[15378] = 210;
razn_w_mem[15379] = 210;
razn_w_mem[15380] = 210;
razn_w_mem[15381] = 210;
razn_w_mem[15382] = 210;
razn_w_mem[15383] = 210;
razn_w_mem[15384] = 210;
razn_w_mem[15385] = 210;
razn_w_mem[15386] = 210;
razn_w_mem[15387] = 210;
razn_w_mem[15388] = 210;
razn_w_mem[15389] = 210;
razn_w_mem[15390] = 210;
razn_w_mem[15391] = 210;
razn_w_mem[15392] = 210;
razn_w_mem[15393] = 210;
razn_w_mem[15394] = 210;
razn_w_mem[15395] = 210;
razn_w_mem[15396] = 210;
razn_w_mem[15397] = 210;
razn_w_mem[15398] = 210;
razn_w_mem[15399] = 210;
razn_w_mem[15400] = 210;
razn_w_mem[15401] = 210;
razn_w_mem[15402] = 210;
razn_w_mem[15403] = 210;
razn_w_mem[15404] = 210;
razn_w_mem[15405] = 210;
razn_w_mem[15406] = 210;
razn_w_mem[15407] = 210;
razn_w_mem[15408] = 210;
razn_w_mem[15409] = 210;
razn_w_mem[15410] = 210;
razn_w_mem[15411] = 210;
razn_w_mem[15412] = 210;
razn_w_mem[15413] = 210;
razn_w_mem[15414] = 210;
razn_w_mem[15415] = 210;
razn_w_mem[15416] = 210;
razn_w_mem[15417] = 210;
razn_w_mem[15418] = 210;
razn_w_mem[15419] = 210;
razn_w_mem[15420] = 210;
razn_w_mem[15421] = 210;
razn_w_mem[15422] = 210;
razn_w_mem[15423] = 210;
razn_w_mem[15424] = 210;
razn_w_mem[15425] = 210;
razn_w_mem[15426] = 210;
razn_w_mem[15427] = 210;
razn_w_mem[15428] = 210;
razn_w_mem[15429] = 210;
razn_w_mem[15430] = 210;
razn_w_mem[15431] = 210;
razn_w_mem[15432] = 210;
razn_w_mem[15433] = 210;
razn_w_mem[15434] = 210;
razn_w_mem[15435] = 210;
razn_w_mem[15436] = 210;
razn_w_mem[15437] = 210;
razn_w_mem[15438] = 210;
razn_w_mem[15439] = 210;
razn_w_mem[15440] = 210;
razn_w_mem[15441] = 210;
razn_w_mem[15442] = 210;
razn_w_mem[15443] = 210;
razn_w_mem[15444] = 210;
razn_w_mem[15445] = 210;
razn_w_mem[15446] = 210;
razn_w_mem[15447] = 210;
razn_w_mem[15448] = 210;
razn_w_mem[15449] = 210;
razn_w_mem[15450] = 210;
razn_w_mem[15451] = 210;
razn_w_mem[15452] = 210;
razn_w_mem[15453] = 210;
razn_w_mem[15454] = 210;
razn_w_mem[15455] = 210;
razn_w_mem[15456] = 210;
razn_w_mem[15457] = 210;
razn_w_mem[15458] = 210;
razn_w_mem[15459] = 210;
razn_w_mem[15460] = 210;
razn_w_mem[15461] = 210;
razn_w_mem[15462] = 210;
razn_w_mem[15463] = 210;
razn_w_mem[15464] = 210;
razn_w_mem[15465] = 210;
razn_w_mem[15466] = 210;
razn_w_mem[15467] = 210;
razn_w_mem[15468] = 210;
razn_w_mem[15469] = 210;
razn_w_mem[15470] = 210;
razn_w_mem[15471] = 210;
razn_w_mem[15472] = 210;
razn_w_mem[15473] = 210;
razn_w_mem[15474] = 210;
razn_w_mem[15475] = 210;
razn_w_mem[15476] = 210;
razn_w_mem[15477] = 210;
razn_w_mem[15478] = 210;
razn_w_mem[15479] = 210;
razn_w_mem[15480] = 210;
razn_w_mem[15481] = 210;
razn_w_mem[15482] = 210;
razn_w_mem[15483] = 210;
razn_w_mem[15484] = 210;
razn_w_mem[15485] = 210;
razn_w_mem[15486] = 210;
razn_w_mem[15487] = 210;
razn_w_mem[15488] = 180;
razn_w_mem[15489] = 180;
razn_w_mem[15490] = 180;
razn_w_mem[15491] = 180;
razn_w_mem[15492] = 180;
razn_w_mem[15493] = 180;
razn_w_mem[15494] = 180;
razn_w_mem[15495] = 180;
razn_w_mem[15496] = 180;
razn_w_mem[15497] = 180;
razn_w_mem[15498] = 180;
razn_w_mem[15499] = 180;
razn_w_mem[15500] = 180;
razn_w_mem[15501] = 180;
razn_w_mem[15502] = 180;
razn_w_mem[15503] = 180;
razn_w_mem[15504] = 180;
razn_w_mem[15505] = 180;
razn_w_mem[15506] = 180;
razn_w_mem[15507] = 180;
razn_w_mem[15508] = 180;
razn_w_mem[15509] = 180;
razn_w_mem[15510] = 180;
razn_w_mem[15511] = 180;
razn_w_mem[15512] = 180;
razn_w_mem[15513] = 180;
razn_w_mem[15514] = 180;
razn_w_mem[15515] = 180;
razn_w_mem[15516] = 180;
razn_w_mem[15517] = 180;
razn_w_mem[15518] = 180;
razn_w_mem[15519] = 180;
razn_w_mem[15520] = 180;
razn_w_mem[15521] = 180;
razn_w_mem[15522] = 180;
razn_w_mem[15523] = 180;
razn_w_mem[15524] = 180;
razn_w_mem[15525] = 180;
razn_w_mem[15526] = 180;
razn_w_mem[15527] = 180;
razn_w_mem[15528] = 180;
razn_w_mem[15529] = 180;
razn_w_mem[15530] = 180;
razn_w_mem[15531] = 180;
razn_w_mem[15532] = 180;
razn_w_mem[15533] = 180;
razn_w_mem[15534] = 180;
razn_w_mem[15535] = 180;
razn_w_mem[15536] = 180;
razn_w_mem[15537] = 180;
razn_w_mem[15538] = 180;
razn_w_mem[15539] = 180;
razn_w_mem[15540] = 180;
razn_w_mem[15541] = 180;
razn_w_mem[15542] = 180;
razn_w_mem[15543] = 180;
razn_w_mem[15544] = 180;
razn_w_mem[15545] = 180;
razn_w_mem[15546] = 180;
razn_w_mem[15547] = 180;
razn_w_mem[15548] = 180;
razn_w_mem[15549] = 180;
razn_w_mem[15550] = 180;
razn_w_mem[15551] = 180;
razn_w_mem[15552] = 180;
razn_w_mem[15553] = 180;
razn_w_mem[15554] = 180;
razn_w_mem[15555] = 180;
razn_w_mem[15556] = 180;
razn_w_mem[15557] = 180;
razn_w_mem[15558] = 180;
razn_w_mem[15559] = 180;
razn_w_mem[15560] = 180;
razn_w_mem[15561] = 180;
razn_w_mem[15562] = 180;
razn_w_mem[15563] = 180;
razn_w_mem[15564] = 180;
razn_w_mem[15565] = 180;
razn_w_mem[15566] = 180;
razn_w_mem[15567] = 180;
razn_w_mem[15568] = 180;
razn_w_mem[15569] = 180;
razn_w_mem[15570] = 180;
razn_w_mem[15571] = 180;
razn_w_mem[15572] = 180;
razn_w_mem[15573] = 180;
razn_w_mem[15574] = 180;
razn_w_mem[15575] = 180;
razn_w_mem[15576] = 180;
razn_w_mem[15577] = 180;
razn_w_mem[15578] = 180;
razn_w_mem[15579] = 180;
razn_w_mem[15580] = 180;
razn_w_mem[15581] = 180;
razn_w_mem[15582] = 180;
razn_w_mem[15583] = 180;
razn_w_mem[15584] = 180;
razn_w_mem[15585] = 180;
razn_w_mem[15586] = 180;
razn_w_mem[15587] = 180;
razn_w_mem[15588] = 180;
razn_w_mem[15589] = 180;
razn_w_mem[15590] = 180;
razn_w_mem[15591] = 180;
razn_w_mem[15592] = 180;
razn_w_mem[15593] = 180;
razn_w_mem[15594] = 180;
razn_w_mem[15595] = 180;
razn_w_mem[15596] = 180;
razn_w_mem[15597] = 180;
razn_w_mem[15598] = 180;
razn_w_mem[15599] = 180;
razn_w_mem[15600] = 180;
razn_w_mem[15601] = 180;
razn_w_mem[15602] = 180;
razn_w_mem[15603] = 180;
razn_w_mem[15604] = 180;
razn_w_mem[15605] = 180;
razn_w_mem[15606] = 180;
razn_w_mem[15607] = 180;
razn_w_mem[15608] = 180;
razn_w_mem[15609] = 180;
razn_w_mem[15610] = 180;
razn_w_mem[15611] = 180;
razn_w_mem[15612] = 180;
razn_w_mem[15613] = 180;
razn_w_mem[15614] = 180;
razn_w_mem[15615] = 180;
razn_w_mem[15616] = 150;
razn_w_mem[15617] = 150;
razn_w_mem[15618] = 150;
razn_w_mem[15619] = 150;
razn_w_mem[15620] = 150;
razn_w_mem[15621] = 150;
razn_w_mem[15622] = 150;
razn_w_mem[15623] = 150;
razn_w_mem[15624] = 150;
razn_w_mem[15625] = 150;
razn_w_mem[15626] = 150;
razn_w_mem[15627] = 150;
razn_w_mem[15628] = 150;
razn_w_mem[15629] = 150;
razn_w_mem[15630] = 150;
razn_w_mem[15631] = 150;
razn_w_mem[15632] = 150;
razn_w_mem[15633] = 150;
razn_w_mem[15634] = 150;
razn_w_mem[15635] = 150;
razn_w_mem[15636] = 150;
razn_w_mem[15637] = 150;
razn_w_mem[15638] = 150;
razn_w_mem[15639] = 150;
razn_w_mem[15640] = 150;
razn_w_mem[15641] = 150;
razn_w_mem[15642] = 150;
razn_w_mem[15643] = 150;
razn_w_mem[15644] = 150;
razn_w_mem[15645] = 150;
razn_w_mem[15646] = 150;
razn_w_mem[15647] = 150;
razn_w_mem[15648] = 150;
razn_w_mem[15649] = 150;
razn_w_mem[15650] = 150;
razn_w_mem[15651] = 150;
razn_w_mem[15652] = 150;
razn_w_mem[15653] = 150;
razn_w_mem[15654] = 150;
razn_w_mem[15655] = 150;
razn_w_mem[15656] = 150;
razn_w_mem[15657] = 150;
razn_w_mem[15658] = 150;
razn_w_mem[15659] = 150;
razn_w_mem[15660] = 150;
razn_w_mem[15661] = 150;
razn_w_mem[15662] = 150;
razn_w_mem[15663] = 150;
razn_w_mem[15664] = 150;
razn_w_mem[15665] = 150;
razn_w_mem[15666] = 150;
razn_w_mem[15667] = 150;
razn_w_mem[15668] = 150;
razn_w_mem[15669] = 150;
razn_w_mem[15670] = 150;
razn_w_mem[15671] = 150;
razn_w_mem[15672] = 150;
razn_w_mem[15673] = 150;
razn_w_mem[15674] = 150;
razn_w_mem[15675] = 150;
razn_w_mem[15676] = 150;
razn_w_mem[15677] = 150;
razn_w_mem[15678] = 150;
razn_w_mem[15679] = 150;
razn_w_mem[15680] = 150;
razn_w_mem[15681] = 150;
razn_w_mem[15682] = 150;
razn_w_mem[15683] = 150;
razn_w_mem[15684] = 150;
razn_w_mem[15685] = 150;
razn_w_mem[15686] = 150;
razn_w_mem[15687] = 150;
razn_w_mem[15688] = 150;
razn_w_mem[15689] = 150;
razn_w_mem[15690] = 150;
razn_w_mem[15691] = 150;
razn_w_mem[15692] = 150;
razn_w_mem[15693] = 150;
razn_w_mem[15694] = 150;
razn_w_mem[15695] = 150;
razn_w_mem[15696] = 150;
razn_w_mem[15697] = 150;
razn_w_mem[15698] = 150;
razn_w_mem[15699] = 150;
razn_w_mem[15700] = 150;
razn_w_mem[15701] = 150;
razn_w_mem[15702] = 150;
razn_w_mem[15703] = 150;
razn_w_mem[15704] = 150;
razn_w_mem[15705] = 150;
razn_w_mem[15706] = 150;
razn_w_mem[15707] = 150;
razn_w_mem[15708] = 150;
razn_w_mem[15709] = 150;
razn_w_mem[15710] = 150;
razn_w_mem[15711] = 150;
razn_w_mem[15712] = 150;
razn_w_mem[15713] = 150;
razn_w_mem[15714] = 150;
razn_w_mem[15715] = 150;
razn_w_mem[15716] = 150;
razn_w_mem[15717] = 150;
razn_w_mem[15718] = 150;
razn_w_mem[15719] = 150;
razn_w_mem[15720] = 150;
razn_w_mem[15721] = 150;
razn_w_mem[15722] = 150;
razn_w_mem[15723] = 150;
razn_w_mem[15724] = 150;
razn_w_mem[15725] = 150;
razn_w_mem[15726] = 150;
razn_w_mem[15727] = 150;
razn_w_mem[15728] = 150;
razn_w_mem[15729] = 150;
razn_w_mem[15730] = 150;
razn_w_mem[15731] = 150;
razn_w_mem[15732] = 150;
razn_w_mem[15733] = 150;
razn_w_mem[15734] = 150;
razn_w_mem[15735] = 150;
razn_w_mem[15736] = 150;
razn_w_mem[15737] = 150;
razn_w_mem[15738] = 150;
razn_w_mem[15739] = 150;
razn_w_mem[15740] = 150;
razn_w_mem[15741] = 150;
razn_w_mem[15742] = 150;
razn_w_mem[15743] = 150;
razn_w_mem[15744] = 120;
razn_w_mem[15745] = 120;
razn_w_mem[15746] = 120;
razn_w_mem[15747] = 120;
razn_w_mem[15748] = 120;
razn_w_mem[15749] = 120;
razn_w_mem[15750] = 120;
razn_w_mem[15751] = 120;
razn_w_mem[15752] = 120;
razn_w_mem[15753] = 120;
razn_w_mem[15754] = 120;
razn_w_mem[15755] = 120;
razn_w_mem[15756] = 120;
razn_w_mem[15757] = 120;
razn_w_mem[15758] = 120;
razn_w_mem[15759] = 120;
razn_w_mem[15760] = 120;
razn_w_mem[15761] = 120;
razn_w_mem[15762] = 120;
razn_w_mem[15763] = 120;
razn_w_mem[15764] = 120;
razn_w_mem[15765] = 120;
razn_w_mem[15766] = 120;
razn_w_mem[15767] = 120;
razn_w_mem[15768] = 120;
razn_w_mem[15769] = 120;
razn_w_mem[15770] = 120;
razn_w_mem[15771] = 120;
razn_w_mem[15772] = 120;
razn_w_mem[15773] = 120;
razn_w_mem[15774] = 120;
razn_w_mem[15775] = 120;
razn_w_mem[15776] = 120;
razn_w_mem[15777] = 120;
razn_w_mem[15778] = 120;
razn_w_mem[15779] = 120;
razn_w_mem[15780] = 120;
razn_w_mem[15781] = 120;
razn_w_mem[15782] = 120;
razn_w_mem[15783] = 120;
razn_w_mem[15784] = 120;
razn_w_mem[15785] = 120;
razn_w_mem[15786] = 120;
razn_w_mem[15787] = 120;
razn_w_mem[15788] = 120;
razn_w_mem[15789] = 120;
razn_w_mem[15790] = 120;
razn_w_mem[15791] = 120;
razn_w_mem[15792] = 120;
razn_w_mem[15793] = 120;
razn_w_mem[15794] = 120;
razn_w_mem[15795] = 120;
razn_w_mem[15796] = 120;
razn_w_mem[15797] = 120;
razn_w_mem[15798] = 120;
razn_w_mem[15799] = 120;
razn_w_mem[15800] = 120;
razn_w_mem[15801] = 120;
razn_w_mem[15802] = 120;
razn_w_mem[15803] = 120;
razn_w_mem[15804] = 120;
razn_w_mem[15805] = 120;
razn_w_mem[15806] = 120;
razn_w_mem[15807] = 120;
razn_w_mem[15808] = 120;
razn_w_mem[15809] = 120;
razn_w_mem[15810] = 120;
razn_w_mem[15811] = 120;
razn_w_mem[15812] = 120;
razn_w_mem[15813] = 120;
razn_w_mem[15814] = 120;
razn_w_mem[15815] = 120;
razn_w_mem[15816] = 120;
razn_w_mem[15817] = 120;
razn_w_mem[15818] = 120;
razn_w_mem[15819] = 120;
razn_w_mem[15820] = 120;
razn_w_mem[15821] = 120;
razn_w_mem[15822] = 120;
razn_w_mem[15823] = 120;
razn_w_mem[15824] = 120;
razn_w_mem[15825] = 120;
razn_w_mem[15826] = 120;
razn_w_mem[15827] = 120;
razn_w_mem[15828] = 120;
razn_w_mem[15829] = 120;
razn_w_mem[15830] = 120;
razn_w_mem[15831] = 120;
razn_w_mem[15832] = 120;
razn_w_mem[15833] = 120;
razn_w_mem[15834] = 120;
razn_w_mem[15835] = 120;
razn_w_mem[15836] = 120;
razn_w_mem[15837] = 120;
razn_w_mem[15838] = 120;
razn_w_mem[15839] = 120;
razn_w_mem[15840] = 120;
razn_w_mem[15841] = 120;
razn_w_mem[15842] = 120;
razn_w_mem[15843] = 120;
razn_w_mem[15844] = 120;
razn_w_mem[15845] = 120;
razn_w_mem[15846] = 120;
razn_w_mem[15847] = 120;
razn_w_mem[15848] = 120;
razn_w_mem[15849] = 120;
razn_w_mem[15850] = 120;
razn_w_mem[15851] = 120;
razn_w_mem[15852] = 120;
razn_w_mem[15853] = 120;
razn_w_mem[15854] = 120;
razn_w_mem[15855] = 120;
razn_w_mem[15856] = 120;
razn_w_mem[15857] = 120;
razn_w_mem[15858] = 120;
razn_w_mem[15859] = 120;
razn_w_mem[15860] = 120;
razn_w_mem[15861] = 120;
razn_w_mem[15862] = 120;
razn_w_mem[15863] = 120;
razn_w_mem[15864] = 120;
razn_w_mem[15865] = 120;
razn_w_mem[15866] = 120;
razn_w_mem[15867] = 120;
razn_w_mem[15868] = 120;
razn_w_mem[15869] = 120;
razn_w_mem[15870] = 120;
razn_w_mem[15871] = 120;
razn_w_mem[15872] = 90;
razn_w_mem[15873] = 90;
razn_w_mem[15874] = 90;
razn_w_mem[15875] = 90;
razn_w_mem[15876] = 90;
razn_w_mem[15877] = 90;
razn_w_mem[15878] = 90;
razn_w_mem[15879] = 90;
razn_w_mem[15880] = 90;
razn_w_mem[15881] = 90;
razn_w_mem[15882] = 90;
razn_w_mem[15883] = 90;
razn_w_mem[15884] = 90;
razn_w_mem[15885] = 90;
razn_w_mem[15886] = 90;
razn_w_mem[15887] = 90;
razn_w_mem[15888] = 90;
razn_w_mem[15889] = 90;
razn_w_mem[15890] = 90;
razn_w_mem[15891] = 90;
razn_w_mem[15892] = 90;
razn_w_mem[15893] = 90;
razn_w_mem[15894] = 90;
razn_w_mem[15895] = 90;
razn_w_mem[15896] = 90;
razn_w_mem[15897] = 90;
razn_w_mem[15898] = 90;
razn_w_mem[15899] = 90;
razn_w_mem[15900] = 90;
razn_w_mem[15901] = 90;
razn_w_mem[15902] = 90;
razn_w_mem[15903] = 90;
razn_w_mem[15904] = 90;
razn_w_mem[15905] = 90;
razn_w_mem[15906] = 90;
razn_w_mem[15907] = 90;
razn_w_mem[15908] = 90;
razn_w_mem[15909] = 90;
razn_w_mem[15910] = 90;
razn_w_mem[15911] = 90;
razn_w_mem[15912] = 90;
razn_w_mem[15913] = 90;
razn_w_mem[15914] = 90;
razn_w_mem[15915] = 90;
razn_w_mem[15916] = 90;
razn_w_mem[15917] = 90;
razn_w_mem[15918] = 90;
razn_w_mem[15919] = 90;
razn_w_mem[15920] = 90;
razn_w_mem[15921] = 90;
razn_w_mem[15922] = 90;
razn_w_mem[15923] = 90;
razn_w_mem[15924] = 90;
razn_w_mem[15925] = 90;
razn_w_mem[15926] = 90;
razn_w_mem[15927] = 90;
razn_w_mem[15928] = 90;
razn_w_mem[15929] = 90;
razn_w_mem[15930] = 90;
razn_w_mem[15931] = 90;
razn_w_mem[15932] = 90;
razn_w_mem[15933] = 90;
razn_w_mem[15934] = 90;
razn_w_mem[15935] = 90;
razn_w_mem[15936] = 90;
razn_w_mem[15937] = 90;
razn_w_mem[15938] = 90;
razn_w_mem[15939] = 90;
razn_w_mem[15940] = 90;
razn_w_mem[15941] = 90;
razn_w_mem[15942] = 90;
razn_w_mem[15943] = 90;
razn_w_mem[15944] = 90;
razn_w_mem[15945] = 90;
razn_w_mem[15946] = 90;
razn_w_mem[15947] = 90;
razn_w_mem[15948] = 90;
razn_w_mem[15949] = 90;
razn_w_mem[15950] = 90;
razn_w_mem[15951] = 90;
razn_w_mem[15952] = 90;
razn_w_mem[15953] = 90;
razn_w_mem[15954] = 90;
razn_w_mem[15955] = 90;
razn_w_mem[15956] = 90;
razn_w_mem[15957] = 90;
razn_w_mem[15958] = 90;
razn_w_mem[15959] = 90;
razn_w_mem[15960] = 90;
razn_w_mem[15961] = 90;
razn_w_mem[15962] = 90;
razn_w_mem[15963] = 90;
razn_w_mem[15964] = 90;
razn_w_mem[15965] = 90;
razn_w_mem[15966] = 90;
razn_w_mem[15967] = 90;
razn_w_mem[15968] = 90;
razn_w_mem[15969] = 90;
razn_w_mem[15970] = 90;
razn_w_mem[15971] = 90;
razn_w_mem[15972] = 90;
razn_w_mem[15973] = 90;
razn_w_mem[15974] = 90;
razn_w_mem[15975] = 90;
razn_w_mem[15976] = 90;
razn_w_mem[15977] = 90;
razn_w_mem[15978] = 90;
razn_w_mem[15979] = 90;
razn_w_mem[15980] = 90;
razn_w_mem[15981] = 90;
razn_w_mem[15982] = 90;
razn_w_mem[15983] = 90;
razn_w_mem[15984] = 90;
razn_w_mem[15985] = 90;
razn_w_mem[15986] = 90;
razn_w_mem[15987] = 90;
razn_w_mem[15988] = 90;
razn_w_mem[15989] = 90;
razn_w_mem[15990] = 90;
razn_w_mem[15991] = 90;
razn_w_mem[15992] = 90;
razn_w_mem[15993] = 90;
razn_w_mem[15994] = 90;
razn_w_mem[15995] = 90;
razn_w_mem[15996] = 90;
razn_w_mem[15997] = 90;
razn_w_mem[15998] = 90;
razn_w_mem[15999] = 90;
razn_w_mem[16000] = 60;
razn_w_mem[16001] = 60;
razn_w_mem[16002] = 60;
razn_w_mem[16003] = 60;
razn_w_mem[16004] = 60;
razn_w_mem[16005] = 60;
razn_w_mem[16006] = 60;
razn_w_mem[16007] = 60;
razn_w_mem[16008] = 60;
razn_w_mem[16009] = 60;
razn_w_mem[16010] = 60;
razn_w_mem[16011] = 60;
razn_w_mem[16012] = 60;
razn_w_mem[16013] = 60;
razn_w_mem[16014] = 60;
razn_w_mem[16015] = 60;
razn_w_mem[16016] = 60;
razn_w_mem[16017] = 60;
razn_w_mem[16018] = 60;
razn_w_mem[16019] = 60;
razn_w_mem[16020] = 60;
razn_w_mem[16021] = 60;
razn_w_mem[16022] = 60;
razn_w_mem[16023] = 60;
razn_w_mem[16024] = 60;
razn_w_mem[16025] = 60;
razn_w_mem[16026] = 60;
razn_w_mem[16027] = 60;
razn_w_mem[16028] = 60;
razn_w_mem[16029] = 60;
razn_w_mem[16030] = 60;
razn_w_mem[16031] = 60;
razn_w_mem[16032] = 60;
razn_w_mem[16033] = 60;
razn_w_mem[16034] = 60;
razn_w_mem[16035] = 60;
razn_w_mem[16036] = 60;
razn_w_mem[16037] = 60;
razn_w_mem[16038] = 60;
razn_w_mem[16039] = 60;
razn_w_mem[16040] = 60;
razn_w_mem[16041] = 60;
razn_w_mem[16042] = 60;
razn_w_mem[16043] = 60;
razn_w_mem[16044] = 60;
razn_w_mem[16045] = 60;
razn_w_mem[16046] = 60;
razn_w_mem[16047] = 60;
razn_w_mem[16048] = 60;
razn_w_mem[16049] = 60;
razn_w_mem[16050] = 60;
razn_w_mem[16051] = 60;
razn_w_mem[16052] = 60;
razn_w_mem[16053] = 60;
razn_w_mem[16054] = 60;
razn_w_mem[16055] = 60;
razn_w_mem[16056] = 60;
razn_w_mem[16057] = 60;
razn_w_mem[16058] = 60;
razn_w_mem[16059] = 60;
razn_w_mem[16060] = 60;
razn_w_mem[16061] = 60;
razn_w_mem[16062] = 60;
razn_w_mem[16063] = 60;
razn_w_mem[16064] = 60;
razn_w_mem[16065] = 60;
razn_w_mem[16066] = 60;
razn_w_mem[16067] = 60;
razn_w_mem[16068] = 60;
razn_w_mem[16069] = 60;
razn_w_mem[16070] = 60;
razn_w_mem[16071] = 60;
razn_w_mem[16072] = 60;
razn_w_mem[16073] = 60;
razn_w_mem[16074] = 60;
razn_w_mem[16075] = 60;
razn_w_mem[16076] = 60;
razn_w_mem[16077] = 60;
razn_w_mem[16078] = 60;
razn_w_mem[16079] = 60;
razn_w_mem[16080] = 60;
razn_w_mem[16081] = 60;
razn_w_mem[16082] = 60;
razn_w_mem[16083] = 60;
razn_w_mem[16084] = 60;
razn_w_mem[16085] = 60;
razn_w_mem[16086] = 60;
razn_w_mem[16087] = 60;
razn_w_mem[16088] = 60;
razn_w_mem[16089] = 60;
razn_w_mem[16090] = 60;
razn_w_mem[16091] = 60;
razn_w_mem[16092] = 60;
razn_w_mem[16093] = 60;
razn_w_mem[16094] = 60;
razn_w_mem[16095] = 60;
razn_w_mem[16096] = 60;
razn_w_mem[16097] = 60;
razn_w_mem[16098] = 60;
razn_w_mem[16099] = 60;
razn_w_mem[16100] = 60;
razn_w_mem[16101] = 60;
razn_w_mem[16102] = 60;
razn_w_mem[16103] = 60;
razn_w_mem[16104] = 60;
razn_w_mem[16105] = 60;
razn_w_mem[16106] = 60;
razn_w_mem[16107] = 60;
razn_w_mem[16108] = 60;
razn_w_mem[16109] = 60;
razn_w_mem[16110] = 60;
razn_w_mem[16111] = 60;
razn_w_mem[16112] = 60;
razn_w_mem[16113] = 60;
razn_w_mem[16114] = 60;
razn_w_mem[16115] = 60;
razn_w_mem[16116] = 60;
razn_w_mem[16117] = 60;
razn_w_mem[16118] = 60;
razn_w_mem[16119] = 60;
razn_w_mem[16120] = 60;
razn_w_mem[16121] = 60;
razn_w_mem[16122] = 60;
razn_w_mem[16123] = 60;
razn_w_mem[16124] = 60;
razn_w_mem[16125] = 60;
razn_w_mem[16126] = 60;
razn_w_mem[16127] = 60;
razn_w_mem[16128] = 30;
razn_w_mem[16129] = 30;
razn_w_mem[16130] = 30;
razn_w_mem[16131] = 30;
razn_w_mem[16132] = 30;
razn_w_mem[16133] = 30;
razn_w_mem[16134] = 30;
razn_w_mem[16135] = 30;
razn_w_mem[16136] = 30;
razn_w_mem[16137] = 30;
razn_w_mem[16138] = 30;
razn_w_mem[16139] = 30;
razn_w_mem[16140] = 30;
razn_w_mem[16141] = 30;
razn_w_mem[16142] = 30;
razn_w_mem[16143] = 30;
razn_w_mem[16144] = 30;
razn_w_mem[16145] = 30;
razn_w_mem[16146] = 30;
razn_w_mem[16147] = 30;
razn_w_mem[16148] = 30;
razn_w_mem[16149] = 30;
razn_w_mem[16150] = 30;
razn_w_mem[16151] = 30;
razn_w_mem[16152] = 30;
razn_w_mem[16153] = 30;
razn_w_mem[16154] = 30;
razn_w_mem[16155] = 30;
razn_w_mem[16156] = 30;
razn_w_mem[16157] = 30;
razn_w_mem[16158] = 30;
razn_w_mem[16159] = 30;
razn_w_mem[16160] = 30;
razn_w_mem[16161] = 30;
razn_w_mem[16162] = 30;
razn_w_mem[16163] = 30;
razn_w_mem[16164] = 30;
razn_w_mem[16165] = 30;
razn_w_mem[16166] = 30;
razn_w_mem[16167] = 30;
razn_w_mem[16168] = 30;
razn_w_mem[16169] = 30;
razn_w_mem[16170] = 30;
razn_w_mem[16171] = 30;
razn_w_mem[16172] = 30;
razn_w_mem[16173] = 30;
razn_w_mem[16174] = 30;
razn_w_mem[16175] = 30;
razn_w_mem[16176] = 30;
razn_w_mem[16177] = 30;
razn_w_mem[16178] = 30;
razn_w_mem[16179] = 30;
razn_w_mem[16180] = 30;
razn_w_mem[16181] = 30;
razn_w_mem[16182] = 30;
razn_w_mem[16183] = 30;
razn_w_mem[16184] = 30;
razn_w_mem[16185] = 30;
razn_w_mem[16186] = 30;
razn_w_mem[16187] = 30;
razn_w_mem[16188] = 30;
razn_w_mem[16189] = 30;
razn_w_mem[16190] = 30;
razn_w_mem[16191] = 30;
razn_w_mem[16192] = 30;
razn_w_mem[16193] = 30;
razn_w_mem[16194] = 30;
razn_w_mem[16195] = 30;
razn_w_mem[16196] = 30;
razn_w_mem[16197] = 30;
razn_w_mem[16198] = 30;
razn_w_mem[16199] = 30;
razn_w_mem[16200] = 30;
razn_w_mem[16201] = 30;
razn_w_mem[16202] = 30;
razn_w_mem[16203] = 30;
razn_w_mem[16204] = 30;
razn_w_mem[16205] = 30;
razn_w_mem[16206] = 30;
razn_w_mem[16207] = 30;
razn_w_mem[16208] = 30;
razn_w_mem[16209] = 30;
razn_w_mem[16210] = 30;
razn_w_mem[16211] = 30;
razn_w_mem[16212] = 30;
razn_w_mem[16213] = 30;
razn_w_mem[16214] = 30;
razn_w_mem[16215] = 30;
razn_w_mem[16216] = 30;
razn_w_mem[16217] = 30;
razn_w_mem[16218] = 30;
razn_w_mem[16219] = 30;
razn_w_mem[16220] = 30;
razn_w_mem[16221] = 30;
razn_w_mem[16222] = 30;
razn_w_mem[16223] = 30;
razn_w_mem[16224] = 30;
razn_w_mem[16225] = 30;
razn_w_mem[16226] = 30;
razn_w_mem[16227] = 30;
razn_w_mem[16228] = 30;
razn_w_mem[16229] = 30;
razn_w_mem[16230] = 30;
razn_w_mem[16231] = 30;
razn_w_mem[16232] = 30;
razn_w_mem[16233] = 30;
razn_w_mem[16234] = 30;
razn_w_mem[16235] = 30;
razn_w_mem[16236] = 30;
razn_w_mem[16237] = 30;
razn_w_mem[16238] = 30;
razn_w_mem[16239] = 30;
razn_w_mem[16240] = 30;
razn_w_mem[16241] = 30;
razn_w_mem[16242] = 30;
razn_w_mem[16243] = 30;
razn_w_mem[16244] = 30;
razn_w_mem[16245] = 30;
razn_w_mem[16246] = 30;
razn_w_mem[16247] = 30;
razn_w_mem[16248] = 30;
razn_w_mem[16249] = 30;
razn_w_mem[16250] = 30;
razn_w_mem[16251] = 30;
razn_w_mem[16252] = 30;
razn_w_mem[16253] = 30;
razn_w_mem[16254] = 30;
razn_w_mem[16255] = 30;
razn_w_mem[16256] = 255;
razn_w_mem[16257] = 255;
razn_w_mem[16258] = 255;
razn_w_mem[16259] = 255;
razn_w_mem[16260] = 255;
razn_w_mem[16261] = 255;
razn_w_mem[16262] = 255;
razn_w_mem[16263] = 255;
razn_w_mem[16264] = 255;
razn_w_mem[16265] = 255;
razn_w_mem[16266] = 255;
razn_w_mem[16267] = 255;
razn_w_mem[16268] = 255;
razn_w_mem[16269] = 255;
razn_w_mem[16270] = 255;
razn_w_mem[16271] = 255;
razn_w_mem[16272] = 255;
razn_w_mem[16273] = 255;
razn_w_mem[16274] = 255;
razn_w_mem[16275] = 255;
razn_w_mem[16276] = 255;
razn_w_mem[16277] = 255;
razn_w_mem[16278] = 255;
razn_w_mem[16279] = 255;
razn_w_mem[16280] = 255;
razn_w_mem[16281] = 255;
razn_w_mem[16282] = 255;
razn_w_mem[16283] = 255;
razn_w_mem[16284] = 255;
razn_w_mem[16285] = 255;
razn_w_mem[16286] = 255;
razn_w_mem[16287] = 255;
razn_w_mem[16288] = 255;
razn_w_mem[16289] = 255;
razn_w_mem[16290] = 255;
razn_w_mem[16291] = 255;
razn_w_mem[16292] = 255;
razn_w_mem[16293] = 255;
razn_w_mem[16294] = 255;
razn_w_mem[16295] = 255;
razn_w_mem[16296] = 255;
razn_w_mem[16297] = 255;
razn_w_mem[16298] = 255;
razn_w_mem[16299] = 255;
razn_w_mem[16300] = 255;
razn_w_mem[16301] = 255;
razn_w_mem[16302] = 255;
razn_w_mem[16303] = 255;
razn_w_mem[16304] = 255;
razn_w_mem[16305] = 255;
razn_w_mem[16306] = 255;
razn_w_mem[16307] = 255;
razn_w_mem[16308] = 255;
razn_w_mem[16309] = 255;
razn_w_mem[16310] = 255;
razn_w_mem[16311] = 255;
razn_w_mem[16312] = 255;
razn_w_mem[16313] = 255;
razn_w_mem[16314] = 255;
razn_w_mem[16315] = 255;
razn_w_mem[16316] = 255;
razn_w_mem[16317] = 255;
razn_w_mem[16318] = 255;
razn_w_mem[16319] = 255;
razn_w_mem[16320] = 255;
razn_w_mem[16321] = 255;
razn_w_mem[16322] = 255;
razn_w_mem[16323] = 255;
razn_w_mem[16324] = 255;
razn_w_mem[16325] = 255;
razn_w_mem[16326] = 255;
razn_w_mem[16327] = 255;
razn_w_mem[16328] = 255;
razn_w_mem[16329] = 255;
razn_w_mem[16330] = 255;
razn_w_mem[16331] = 255;
razn_w_mem[16332] = 255;
razn_w_mem[16333] = 255;
razn_w_mem[16334] = 255;
razn_w_mem[16335] = 255;
razn_w_mem[16336] = 255;
razn_w_mem[16337] = 255;
razn_w_mem[16338] = 255;
razn_w_mem[16339] = 255;
razn_w_mem[16340] = 255;
razn_w_mem[16341] = 255;
razn_w_mem[16342] = 255;
razn_w_mem[16343] = 255;
razn_w_mem[16344] = 255;
razn_w_mem[16345] = 255;
razn_w_mem[16346] = 255;
razn_w_mem[16347] = 255;
razn_w_mem[16348] = 255;
razn_w_mem[16349] = 255;
razn_w_mem[16350] = 255;
razn_w_mem[16351] = 255;
razn_w_mem[16352] = 255;
razn_w_mem[16353] = 255;
razn_w_mem[16354] = 255;
razn_w_mem[16355] = 255;
razn_w_mem[16356] = 255;
razn_w_mem[16357] = 255;
razn_w_mem[16358] = 255;
razn_w_mem[16359] = 255;
razn_w_mem[16360] = 255;
razn_w_mem[16361] = 255;
razn_w_mem[16362] = 255;
razn_w_mem[16363] = 255;
razn_w_mem[16364] = 255;
razn_w_mem[16365] = 255;
razn_w_mem[16366] = 255;
razn_w_mem[16367] = 255;
razn_w_mem[16368] = 255;
razn_w_mem[16369] = 255;
razn_w_mem[16370] = 255;
razn_w_mem[16371] = 255;
razn_w_mem[16372] = 255;
razn_w_mem[16373] = 255;
razn_w_mem[16374] = 255;
razn_w_mem[16375] = 255;
razn_w_mem[16376] = 255;
razn_w_mem[16377] = 255;
razn_w_mem[16378] = 255;
razn_w_mem[16379] = 255;
razn_w_mem[16380] = 255;
razn_w_mem[16381] = 255;
razn_w_mem[16382] = 255;
razn_w_mem[16383] = 255;
end

endmodule