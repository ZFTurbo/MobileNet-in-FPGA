module  ov5640_cfg(
        
);



endmodule